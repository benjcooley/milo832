`timescale 1ns/1ps


`include "../Memory/fifo.sv"

//=============================================================================
// Module: streaming_multiprocessor
//=============================================================================
// Architecture: Advanced 5-stage SIMT GPU Core (Kepler-class)
//
// OVERVIEW:
//   This module implements a sophisticated Streaming Multiprocessor (SM) designed 
//   for high-throughput GPGPU workloads. It executes 32-thread warps in lockstep 
//   using a Single-Instruction, Multiple-Thread (SIMT) model. The architecture 
//   mimics the NVIDIA Kepler/Fermi evolution, featuring dual-issue superscalar 
//   execution, a decoupled operand collector, and asynchronous memory handling.
//
// ARCHITECTURAL SPECIFICATIONS & MECHANISMS:
//
//   1. DUAL-ISSUE WARP SCHEDULER:
//      - Employs a Loose Round-Robin selection policy among ready warps.
//      - Fetches two contiguous 64-bit instructions for the selected warp.
//      - Performs structural hazard detection (port disjointness) and scoreboard 
//        validation to attempt concurrent issue to ALU, LSU, or SFU/FPU backends.
//
//   2. SOPHISTICATED HAZARD MANAGEMENT (Scoreboard):
//      - Implements a precise per-warp Scoreboard tracking all pending register 
//        writes (WAW/RAW protection).
//      - Tracks dependencies across both synchronous (ALU) and asynchronous 
//        (LSU/FPU) pipelines, ensuring strict program order for data dependencies.
//
//   3. FERMI-STYLE OPERAND COLLECTOR (OC):
//      - Decentralizes the Register File (RF) bandwidth bottleneck using 16 
//        shared Collector Units (CUs).
//      - Interleaves the RF into 4 physical banks (Interleaved Banking).
//      - CUs arbitrate for bank access over multiple cycles to assemble a 
//        complete three-operand instruction bundle (rs1, rs2, rs3) before 
//        releasing it to the execution units.
//
//   4. SPECIAL FUNCTION UNIT (SFU) & FPU:
//      - Supports IEEE-754 single-precision floating-point arithmetic (FADD, FMUL, FFMA).
//      - Dedicated SFU lanes provide high-throughput transcendental operations 
//        (SIN, COS, RCP, RSQ, TANH, LG2, EX2).
//      - Math logic utilizes 1.15 fixed-point ROM lookups with hardware-accelerated 
//        linear interpolation and correct sign-extension for 32-bit registers.
//
//   5. SIMT CONTROL FLOW & DIVERGENCE:
//      - Implements the SSY/JOIN convergence model using a per-warp hardware stack.
//      - Automatically manages thread masks during branch divergence, pushing 
//        the "not-taken" path to the stack for later execution.
//      - Features a Hardware Return Address Stack (RAS) for efficient CALL/RET.
//
//   6. NON-BLOCKING MEMORY SUBSYSTEM (MSHR):
//      - Features a non-blocking interface to a mock L1 cache/DRAM system.
//      - Utilizes Miss Status Holding Registers (MSHR) to track up to 64 outstanding 
//        memory transactions per warp.
//      - Supports split-transaction writebacks, allowing other warps to progress 
//        while memory requests are in flight.
//
// PIPELINE TOPOLOGY:
//   [IF] Fetch & Dual-Issue Check -> [ID] Decode & Scoreboard Reserve -> 
//   [OC] Operand Collection & Arbitration -> [EX] Compute/LSU Execute -> 
//   [WB] Asynchronous Writeback & Scoreboard Clear
//=============================================================================
import simt_pkg::*;
import sfu_pkg::*;

module streaming_multiprocessor
#(
    parameter WARP_SIZE = 32,
    parameter NUM_WARPS = 24,
    parameter NUM_REGS = 64,
    parameter DIVERGENCE_STACK_DEPTH = 32,
    parameter RETURN_STACK_DEPTH = 8,
    parameter ADDR_WIDTH = 10,
    parameter MAX_PENDING_PER_WARP = 64,
    parameter SM_ID = 0,
    parameter NUM_COLLECTORS = 32
)(
    input  logic clk,
    input  logic rst_n,
    output logic done
);

    // Derived parameters
    localparam WARP_ID_WIDTH = $clog2(NUM_WARPS);
    localparam REG_ADDR_WIDTH = $clog2(NUM_REGS);
    
    // TX ID Layout Parameters
    localparam SLOT_ID_WIDTH = $clog2(MAX_PENDING_PER_WARP);
    localparam WARP_ID_OFFSET = SLOT_ID_WIDTH; // Slot occupies lowest bits
    localparam SM_ID_OFFSET = WARP_ID_OFFSET + WARP_ID_WIDTH; // Warp ID above Slot ID
    
    // Ensure TX ID fits (16 bits)
    initial begin
        if (SM_ID_OFFSET + 4 > 16) $error("TX ID width exceeded! Reduce parameters.");
    end

    int cycle;
    logic done_prev;

    // Architectural State
    
    // Predicate Registers: 7 predicates per thread (P0-P6). P7 is constant True.
    logic [6:0]  preds [NUM_WARPS][WARP_SIZE];
    
    initial begin
        for(int w=0; w<NUM_WARPS; w++) begin
             for(int l=0; l<WARP_SIZE; l++) preds[w][l] = 0;
        end
    end
    
    // Warp State
    logic [31:0]              warp_pc           [NUM_WARPS];
    warp_state_e              warp_state        [NUM_WARPS];
    logic [WARP_SIZE-1:0]     warp_active_mask  [NUM_WARPS];
    logic [NUM_REGS-1:0]      warp_reg_writes   [NUM_WARPS];
    logic [7:0]               warp_pred_writes  [NUM_WARPS]; // PREDICATE SCOREBOARD
    logic [$clog2(DIVERGENCE_STACK_DEPTH):0] warp_stack_ptr [NUM_WARPS];
    logic [$clog2(RETURN_STACK_DEPTH):0]     warp_ret_ptr   [NUM_WARPS];
    logic                     warp_at_barrier   [NUM_WARPS];
    
    // Branch Tag for Flush Handling
    logic [1:0] warp_branch_tag [NUM_WARPS];
    
    // Stability & Single-Writer Signals
    warp_state_e warp_state_next [NUM_WARPS];
    logic        init_phase;
    logic        done_next;
    
    logic [NUM_WARPS-1:0] state_req_exit;
    logic [NUM_WARPS-1:0] state_req_barrier;
    logic [NUM_WARPS-1:0] state_req_ready;
    
    // Registered stabilization signals
    logic [NUM_WARPS-1:0][NUM_REGS-1:0] reg_clear_q;
    logic [1:0]                         oc_wb_valid_q;
    logic [1:0][WARP_ID_WIDTH-1:0]      oc_wb_warp_q;
    logic [1:0][REG_ADDR_WIDTH-1:0]     oc_wb_rd_q;
    logic [1:0][WARP_SIZE-1:0]          oc_wb_mask_q;
    logic [1:0][WARP_SIZE-1:0][31:0]    oc_wb_result_q;
    logic [1:0]                         oc_wb_we_q;
    logic [1:0]                         oc_wb_we_pred_q;
    
    
    logic [31:0]          stack_pc   [NUM_WARPS][DIVERGENCE_STACK_DEPTH];
    logic [WARP_SIZE-1:0] stack_mask [NUM_WARPS][DIVERGENCE_STACK_DEPTH];
    logic [31:0]          ret_stack  [NUM_WARPS][RETURN_STACK_DEPTH];  // Return address stack for CALL/RET
    
    
    // Signals for Async Writeback Scoreboard Update
    logic       async_wb_en;
    logic [4:0] async_wb_warp;
    logic [7:0] async_wb_rd;
    
    // MSHR: Fixed Size Table per Warp (Avoids Verilator dynamic queue bug)
    // Indexed by Slot ID (TxID lowest bits)
    pending_load_t mshr_table [NUM_WARPS][MAX_PENDING_PER_WARP]; 
    logic [MAX_PENDING_PER_WARP-1:0] mshr_valid [NUM_WARPS];
    int mshr_count [NUM_WARPS];
    
    // TX ID FIFO Signals
    localparam TX_ID_WIDTH = 16;
    logic [TX_ID_WIDTH-1:0] tx_id_fifo_din  [NUM_WARPS];
    logic [TX_ID_WIDTH-1:0] tx_id_fifo_dout [NUM_WARPS];
    logic                   tx_id_fifo_push [NUM_WARPS];
    logic                   tx_id_fifo_pop  [NUM_WARPS];
    logic                   tx_id_fifo_full [NUM_WARPS];
    logic                   tx_id_fifo_empty[NUM_WARPS];
    int                     tx_id_fifo_count[NUM_WARPS];
    
    // FIFO Driver Signals (Multiple Sources)
    logic                   alloc_pop      [NUM_WARPS];
    logic                   reclaim_push   [NUM_WARPS];
    logic [TX_ID_WIDTH-1:0] reclaim_data   [NUM_WARPS];
    logic                   init_push      [NUM_WARPS];
    logic [TX_ID_WIDTH-1:0] init_data      [NUM_WARPS];

    // MUX Logic for FIFO Inputs
    always_comb begin
        for (int w=0; w<NUM_WARPS; w++) begin
            // 1. Pop Logic: Allocation pops. 
            // FIXED: Only pop if we are NOT in init phase and not pushing (or handling properly)
            // But wait, the user said arbitrate explicitly.
            tx_id_fifo_pop[w]  = alloc_pop[w];
            
            // 2. Push Logic: Init OR Reclaim
            // PRIORITY: Init Phase > Reclaim (Mutual Exclusion strictly enforced by cycle)
            if (cycle < MAX_PENDING_PER_WARP + 2) begin // Init Phase
                tx_id_fifo_push[w] = init_push[w];
                tx_id_fifo_din[w]  = init_data[w];
            end else begin // Run Phase
                // Reclaim Push Logic
                tx_id_fifo_push[w] = reclaim_push[w];
                tx_id_fifo_din[w]  = reclaim_data[w];
            end
        end
    end

    // Instantiate FIFO per Warp
    generate
        for (genvar w=0; w<NUM_WARPS; w++) begin : gen_tx_fifo
            fifo #(
                .DEPTH(MAX_PENDING_PER_WARP),
                .T(logic [TX_ID_WIDTH-1:0])
            ) tx_id_queue (
                .clk(clk),
                .rst_n(rst_n),
                .push(tx_id_fifo_push[w]),
                .pop(tx_id_fifo_pop[w]),
                .data_in(tx_id_fifo_din[w]),
                .data_out(tx_id_fifo_dout[w]),
                .full(tx_id_fifo_full[w]),
                .empty(tx_id_fifo_empty[w]),
                .count(tx_id_fifo_count[w])
            );
        end
    endgenerate


    // Scoreboard Management consolidated into ID stage logic
    
    // ========================================================================
    // Scoreboard Bypass Logic
    // ========================================================================
    // Combinational bypass: Compute which registers are being cleared THIS cycle
    // This allows scoreboard_ok to see clears before they're registered, solving
    // the NBA race condition where scoreboard clears happen in the NBA region
    logic [NUM_WARPS-1:0][NUM_REGS-1:0] reg_clear_this_cycle;
    logic [NUM_WARPS-1:0][7:0]          pred_clear_this_cycle;
    
    always_comb begin
        reg_clear_this_cycle = '0;
        pred_clear_this_cycle = '0;
        
        // Clear Predicate Scoreboard (From ALU WB)
        if (alu_wb.valid && alu_wb.we_pred) begin
            pred_clear_this_cycle[alu_wb.warp][alu_wb.rd[2:0]] = 1;
        end
        
        // Clear Scoreboard from OC Writeback Ports (Sync & Async)
        for (int k=0; k<2; k++) begin
            if (oc_wb_valid[k]) begin
                // ONLY clear if this is the generic ALU/FPU path (always full) 
                // OR if it's a Memory path and this is the LAST split.
                // Note: oc_wb_last_split is needed here.
                // Assuming logic added via implicit wire connection or we decode src
                // For simplified logic: checks specific to Memory WB logic below
                reg_clear_this_cycle[oc_wb_warp[k]][oc_wb_rd[k]] = 1;

                // Optimization: We could qualify with last_split here if we routed it.
                // For now, let's rely on the upstream (Atomic WB) NOT setting Valid if it shouldn't clear?
                // NO. WB must happen for data.
                // We MUST access `mem_resp_wb.last_split`.
                // Port 1 is driven by mem_resp_wb. 
                if (k == 1 && mem_resp_wb.valid) begin
                    // Override: Only clear if last_split is true
                    reg_clear_this_cycle[oc_wb_warp[k]][oc_wb_rd[k]] = mem_resp_wb.last_split;
                end
            end
        end
    end

    // ========================================================================
    // Memory State
    // ========================================================================
    logic [63:0] prog_mem [NUM_WARPS][256];

    // Pipeline Registers (Dual-Issue with Separate ALU/LSU Pipelines)
    if_id_t  if_id[1:0];
    id_ex_t  id_ex[1:0];
    
    // ALU Pipeline: EX → WB (single cycle)
    alu_wb_t alu_wb;
    
    // LSU Pipeline: ADDR → MEM (multi-cycle, async)
    typedef struct packed {
        logic valid;
        logic [4:0] warp;
        opcode_t op;
        logic [7:0] rd;
        logic [WARP_SIZE-1:0] mask;
        logic [WARP_SIZE-1:0][31:0] addresses;
        logic [WARP_SIZE-1:0][31:0] store_data;
    } lsu_mem_t;
    lsu_mem_t lsu_mem;
    
    // Temporary: Keep ex_mem for compatibility during transition
    ex_mem_t ex_mem;
    
    mem_wb_t mem_wb;  // Keep for compatibility (will be phased out)

    // Branch Feedback (EX -> IF)
    logic       branch_taken_q;
    logic [WARP_ID_WIDTH-1:0] branch_warp_q;
    logic [31:0] branch_target_q;

    // Combinational signals generated in EX
    logic       branch_valid_c;
    logic [7:0] branch_target_c;
    
    // Next-state variables for EX Sequential block (Internal Use)
    // --- Branch Signaling (Intermediate) ---
    logic        cur_branch_taken;
    logic [31:0] cur_branch_target;
    logic [WARP_ID_WIDTH-1:0] cur_branch_warp;

    // --- Operand Collector Integration ---
    logic [1:0] oc_dispatch_valid;
    id_ex_t [1:0] oc_dispatch_inst;
    logic [1:0] oc_dispatch_ready;
    
    logic [1:0] oc_ex_valid;
    id_ex_t [1:0] oc_ex_inst;
    logic [1:0] oc_ex_ready;

    // Dual Writeback Signals
    logic [1:0]                      oc_wb_valid;
    logic [1:0][4:0]                 oc_wb_warp;
    logic [1:0][REG_ADDR_WIDTH-1:0]  oc_wb_rd;
    logic [1:0][WARP_SIZE-1:0]       oc_wb_mask;
    logic [1:0][WARP_SIZE-1:0][31:0] oc_wb_data;

    operand_collector #(
        .WARP_SIZE(WARP_SIZE),
        .NUM_REGS(NUM_REGS),
        .NUM_WARPS(NUM_WARPS),
        .NUM_COLLECTORS(NUM_COLLECTORS)
    ) oc_inst (
        .clk(clk),
        .rst_n(rst_n),
        
        .dispatch_valid(oc_dispatch_valid),
        .dispatch_inst(oc_dispatch_inst),
        .dispatch_ready(oc_dispatch_ready),
        
        .wb_valid(oc_wb_valid_q),
        .wb_warp(oc_wb_warp_q),
        .wb_rd(oc_wb_rd_q),
        .wb_mask(oc_wb_mask_q),
        .wb_data(oc_wb_result_q),
        
        .ex_valid(oc_ex_valid),
        .ex_inst(oc_ex_inst),
        .ex_ready(oc_ex_ready),
        
        .flush_valid(1'b0),
        .flush_warp(5'b0),
        .current_warp_branch_tag(warp_branch_tag)
    );

    // Writeback Port 0 (Sync - ALU)
    // Writeback Port 0 (Sync - ALU)
    // Directly driven by ALU Pipeline Register (alu_wb)
    // Writeback Pipeline Registers
    // alu_wb and lsu_mem are declared in Execution Stage Header (lines 193/205)
    // mem_wb_t alu_wb;     // Path A: Compute (ALU) - ALREADY DECLARED
    // mem_wb_t lsu_mem;    // Path B: Memory Request (LSU) - Bridge - ALREADY DECLARED
    mem_wb_t fpu_wb;     // Path C: FPU/SFU
    mem_wb_t mem_resp_wb;// Path D: Memory Response (Async)
    mem_wb_t mem_resp_wb_next; // Next-state for atomic WB
    
    // Writeback Control Signals
    logic fpu_wb_served;
    logic stall_shared_mem_wb;
    assign stall_fpu_wb = fpu_wb.valid && !fpu_wb_served;

    // CENTRAL WRITEBACK ARBITER (Combinational)
    // Updated to detect and prevent Register File Bank Conflicts
    // logic stall_mem_wb; // MOVED TO MODULE LEVEL for feedback
    
    always_comb begin
        oc_wb_valid = 2'b00;
        oc_wb_warp  = '0;
        oc_wb_rd    = '0;
        oc_wb_mask  = '0;
        oc_wb_data  = '0;
        fpu_wb_served = 0;

        // Port 0: Priority ALU -> FPU
        // Use .valid (not .we) to ensure Scoreboard clears even for squashed/predicated-off ops
        if (alu_wb.valid) begin
            oc_wb_valid[0] = 1;
            oc_wb_warp[0]  = alu_wb.warp;
            oc_wb_rd[0]    = alu_wb.rd[REG_ADDR_WIDTH-1:0];
            oc_wb_mask[0]  = alu_wb.we ? alu_wb.mask : '0; 
            oc_wb_data[0]  = alu_wb.result;
        end else if (fpu_wb.valid) begin
            oc_wb_valid[0] = 1;
            oc_wb_warp[0]  = fpu_wb.warp;
            oc_wb_rd[0]    = fpu_wb.rd[REG_ADDR_WIDTH-1:0];
            oc_wb_mask[0]  = fpu_wb.we ? fpu_wb.mask : '0;
            oc_wb_data[0]  = fpu_wb.result;
            fpu_wb_served  = 1;
        end

        // Port 1: Priority MEM_RESP -> FPU
        if (mem_resp_wb.valid) begin
             oc_wb_valid[1] = 1;
             oc_wb_warp[1]  = mem_resp_wb.warp;
             oc_wb_rd[1]    = mem_resp_wb.rd[REG_ADDR_WIDTH-1:0];
             oc_wb_mask[1]  = mem_resp_wb.we ? mem_resp_wb.mask : '0;
             oc_wb_data[1]  = mem_resp_wb.result;
        end else if (fpu_wb.valid && !fpu_wb_served) begin
             oc_wb_valid[1] = 1;
             oc_wb_warp[1]  = fpu_wb.warp;
             oc_wb_rd[1]    = fpu_wb.rd[REG_ADDR_WIDTH-1:0];
             oc_wb_mask[1]  = fpu_wb.we ? fpu_wb.mask : '0;
             oc_wb_data[1]  = fpu_wb.result;
             fpu_wb_served  = 1;
        end
    end

    // Barrier State
    logic [NUM_WARPS-1:0] barrier_mask;
    logic [NUM_WARPS-1:0] barrier_expected; // Tracks warps participating in the CTA
    
    // Barrier Epoch (toggles each completed barrier)
    logic barrier_epoch;
    // Tracks whether a warp has arrived in the current epoch
    logic [NUM_WARPS-1:0] barrier_seen_epoch;
    // Latch signal to freeze barrier_expected on first arrival
    logic barrier_active;
    // Initialization signal to delay release check by one cycle
    logic barrier_initialized;
    
    //=========================================================================
    // PIPELINE STAGE: IF (Instruction Fetch)
    //=========================================================================
    // - Round-robin warp scheduler selects next ready warp
    // - Fetches instruction from program memory
    // - Advances PC for selected warp
    // - Checks scoreboard to avoid issuing instructions with pending operands
    //=========================================================================
    // Round-Robin Pointer
    int rr_ptr;
    
    // Diagnostic Function: Print blocked registers
    function automatic void scoreboard_diag(input int w, input logic [63:0] inst);
        logic [7:0] rs1, rs2, rd, rs3;
        opcode_t op;
        logic rs1_busy, rs2_busy, rs3_busy, rd_busy;
        
        op  = opcode_t'(inst[63:56]);
        rd  = inst[55:48];
        rs1 = inst[47:40];
        rs2 = inst[39:32];
        rs3 = inst[27:20];
        
        rs1_busy = warp_reg_writes[w][ 6'(rs1) ] && !reg_clear_q[w][ 6'(rs1) ];
        rs2_busy = warp_reg_writes[w][ 6'(rs2) ] && !reg_clear_q[w][ 6'(rs2) ];
        rs3_busy = warp_reg_writes[w][ 6'(rs3) ] && !reg_clear_q[w][ 6'(rs3) ];
        rd_busy = warp_reg_writes[w][ 6'(rd) ] && !reg_clear_q[w][ 6'(rd) ];

    $display("CORE [%0t] SB_DIAG: Warp %0d PC=%h Op=%s RS1(%0d)=%b RS2(%0d)=%b RS3(%0d)=%b RD(%0d)=%b", 
                 $time, w, warp_pc[w], op.name(), rs1, rs1_busy, rs2, rs2_busy, rs3, rs3_busy, rd, rd_busy);
        
        // Match in OC
        for (int i=0; i<NUM_COLLECTORS; i++) begin
            if (oc_inst.collectors[i].state != 0 && oc_inst.collectors[i].inst.warp == 5'(w)) begin
                $display("CORE [%0t] OC_MATCH: Unit %0d Warp %0d PC=%h State=%s RS1_Rdy=%b RS2_Rdy=%b RS3_Rdy=%b Needs=%b",
                         $time, i, w, oc_inst.collectors[i].inst.pc, oc_inst.collectors[i].state.name(), 
                         oc_inst.rs1_ready[i], oc_inst.rs2_ready[i], oc_inst.rs3_ready[i], oc_inst.collectors[i].needed_mask);
            end
        end
    endfunction
    

    // Function: Scoreboard Check
    function automatic logic scoreboard_ok(input int w, input logic [63:0] inst);
        logic [7:0] rs1, rs2, rd, rs3;
        opcode_t op;
        logic rs1_busy, rs2_busy, rs3_busy, rd_busy;
        
        op  = opcode_t'(inst[63:56]);
        rd  = inst[55:48];
        rs1 = inst[47:40];
        rs2 = inst[39:32];
        rs3 = inst[27:20];
        
        scoreboard_ok = 1;
        
        if (op != OP_NOP && op != OP_EXIT) begin
            // 0. Predicate Guard Dependency Check
            logic [3:0] pg;
            pg = inst[31:28]; // Predicate Guard Field
            if (pg[2:0] != 7) begin // If not Always True (P7)
                // Check if the predicate register is being written to
                // Note: We check pred_writes vs pred_clear to handle back-to-back
                if (warp_pred_writes[w][pg[2:0]] && !pred_clear_this_cycle[w][pg[2:0]]) begin
                    scoreboard_ok = 0;
                end
            end

            // 1. Initial Busy Check against Registered Scoreboard Clear
            rs1_busy = warp_reg_writes[w][ 6'(rs1) ] && !reg_clear_q[w][ 6'(rs1) ];
            if (op inside {OP_ADD,OP_SUB,OP_MUL,OP_IMAD,OP_SLT,OP_LDR,OP_STR,OP_BEQ,OP_BNE,
                           OP_FADD,OP_FSUB,OP_FMUL,OP_FDIV,OP_FFMA,
                           OP_SFU_SIN,OP_SFU_COS,OP_SFU_RCP,OP_SFU_RSQ,OP_SFU_SQRT,OP_SFU_EX2,OP_SFU_LG2,
                           OP_ITOF,OP_FTOI,OP_IDIV,OP_IREM,OP_IMIN,OP_IMAX,OP_IABS,
                           OP_FMIN,OP_FMAX,OP_FABS,OP_AND,OP_OR,OP_XOR,OP_NOT,
                           OP_SHL,OP_SHR,OP_SHA,OP_POPC,OP_CLZ,OP_BREV,OP_NEG,OP_FNEG,OP_CNOT,
                           OP_SLE,OP_SEQ,OP_ISETP,OP_FSETP,OP_SELP,OP_TID,OP_MOV,OP_LDS,OP_STS} && rs1_busy) 
                scoreboard_ok = 0;
            
            rs2_busy = warp_reg_writes[w][ 6'(rs2) ] && !reg_clear_q[w][ 6'(rs2) ];
            if (op inside {OP_ADD,OP_SUB,OP_MUL,OP_SLT,OP_STR,OP_BEQ,OP_BNE,
                           OP_FADD,OP_FSUB,OP_FMUL,OP_FDIV,OP_FFMA,
                           OP_IDIV,OP_IREM, OP_IMIN,OP_IMAX, OP_FMIN,OP_FMAX,
                           OP_AND,OP_OR,OP_XOR, OP_SHL,OP_SHR,OP_SHA, OP_SLE,OP_SEQ,OP_ISETP,OP_FSETP,OP_STS} && rs2_busy) 
                scoreboard_ok = 0;
                
            rs3_busy = warp_reg_writes[w][ 6'(rs3) ] && !reg_clear_q[w][ 6'(rs3) ];
            if (op inside {OP_FFMA, OP_IMAD} && rs3_busy) scoreboard_ok = 0;
            
            rd_busy = warp_reg_writes[w][ 6'(rd) ] && !reg_clear_q[w][ 6'(rd) ];
            if (op != OP_STR && op != OP_STS && op != OP_BEQ && op != OP_BNE && op != OP_BRA && op != OP_BAR && rd_busy)
                scoreboard_ok = 0;

            // 2. Lookahead Check: Check against instructions in IF/ID stage (not yet reserved in reg_writes)
            for (int p=0; p<2; p++) begin
                if (if_id[p].valid && if_id[p].warp == w[4:0]) begin
                    logic [7:0] if_rd;
                    opcode_t if_op;
                    if_op = opcode_t'(if_id[p].inst[63:56]);
                    if_rd = if_id[p].inst[55:48];
                    
                    // Does if_id[p] write back?
                    if (if_op inside {OP_ADD,OP_SUB,OP_MUL,OP_IMAD,OP_SLT,OP_LDR,OP_STR,OP_TID,
                                     OP_FADD,OP_FSUB,OP_FMUL,OP_FDIV,OP_FFMA,
                                     OP_SFU_SIN,OP_SFU_COS,OP_SFU_RCP,OP_SFU_RSQ,OP_SFU_SQRT,OP_SFU_EX2,OP_SFU_LG2,
                                     OP_ITOF,OP_FTOI,OP_IDIV,OP_IREM,OP_IMIN,OP_IMAX,OP_IABS,
                                     OP_FMIN,OP_FMAX,OP_FABS,OP_AND,OP_OR,OP_XOR,OP_NOT,
                                     OP_SHL,OP_SHR,OP_SHA,OP_POPC,OP_CLZ,OP_BREV,OP_NEG,OP_FNEG,OP_CNOT,
                                     OP_SLE,OP_SEQ,OP_ISETP,OP_FSETP,OP_SELP,OP_MOV,OP_LDS,OP_STS}) begin
                        if (if_rd == rs1 || if_rd == rs2 || if_rd == rs3 || if_rd == rd) begin
                            scoreboard_ok = 0;
                        end
                    end
                    
                    // Predicate RAW Check: If Lookahead instruction writes a predicate we need
                    if (if_op inside {OP_ISETP, OP_FSETP}) begin
                        logic [2:0] if_pred_rd;
                        if_pred_rd = if_id[p].inst[50:48]; // Predicate Destination
                        
                        // Check if we use it as Guard
                        if (pg[2:0] != 7 && pg[2:0] == if_pred_rd) scoreboard_ok = 0;
                        
                        // Check if we use it as Source (SELP)
                        if (op == OP_SELP && inst[2:0] == if_pred_rd) scoreboard_ok = 0;
                    end
                end
            end
        end
    endfunction

    // Function: Check Dual Issue Eligibility
    function automatic logic can_dual_issue(input logic [63:0] inst_a, input logic [63:0] inst_b);
        opcode_t op_a, op_b;
        unit_type_e type_a, type_b;
        
        op_a = opcode_t'(inst_a[63:56]);
        op_b = opcode_t'(inst_b[63:56]);
        
        type_a = get_unit_type(op_a);
        type_b = get_unit_type(op_b);
        
        // Rule: Must target different execution units (Structural Hazard Check)
        // Exceptions can be made if we have multiple units (e.g., 2 ALUs), but currently we route by Type.
        // ALU and CTRL share the ALU/Branch unit.
        // LSU has its own FIFO.
        // FPU/SFU share the Float unit.
        
        if (type_a == type_b) return 0;
        
        // Additional constraint: Control flow instructions usually force single issue in Kepler
        if (type_a == UNIT_CTRL || type_b == UNIT_CTRL) return 0;
        
        return 1;
    endfunction

    // Scheduler Logic
    logic [NUM_WARPS-1:0] issue_eligible_mask;

    // Loop 1: Wakeup Phase (Parallel Eligibility Check)
    always_comb begin
        for (int w=0; w<NUM_WARPS; w++) begin
            issue_eligible_mask[w] = 0;
            if (warp_state[w] == W_READY) begin
                // Efficiency: Check if warp has TX IDs available if it's about to do a memory op
                // This prevents it from being selected only to stall the whole pipeline.
                logic [63:0] next_inst = prog_mem[w][ warp_pc[w][7:0] ];
                opcode_t op = opcode_t'(next_inst[63:56]);
                logic needs_tx_id = (op == OP_LDR || op == OP_STR);
                logic tx_id_ok = !needs_tx_id || !tx_id_fifo_empty[w];

                if (tx_id_ok && scoreboard_ok(int'(w), next_inst)) begin
                    issue_eligible_mask[w] = 1;
                end
            end
        end
    end

    // ========================================================================
    // Warp Scheduler
    // ========================================================================
    // Scheduler state
    logic [WARP_ID_WIDTH-1:0] last_issued_warp;
    logic                     last_issued_valid;

    // Per-warp backpressure: stall if memory op but no TX ID
    logic [NUM_WARPS-1:0] warp_mem_stall;
    
    always_comb begin
        for (int w=0; w<NUM_WARPS; w++) begin
            // Stall this warp if it has a pending memory op but no TX ID available
            warp_mem_stall[w] = (lsu_mem.valid && (lsu_mem.op == OP_LDR || lsu_mem.op == OP_STR) && 
                                (lsu_mem.warp == w) && tx_id_fifo_empty[w]);
        end
    end

    logic stall_pipeline;
    logic fsm_stall;
    logic mem_pool_full_stall;
    logic shared_mem_stall_cpu; // Stall signal from shared_memory serialization
    assign stall_pipeline = fsm_stall || 
                           (oc_dispatch_valid[0] && !oc_dispatch_ready[0]) || 
                           (oc_dispatch_valid[1] && !oc_dispatch_ready[1]) || 
                           shared_mem_stall_cpu;
    
    always_ff @(posedge clk) begin
        if (!oc_dispatch_ready[0] && !rst_n) begin
        end else if (!oc_dispatch_ready[0]) begin
            if (cycle % 100 == 0) $display("CORE [%0t] OC FULL STALL", $time);
        end
    end
    
    // mem_pool_full_stall is now handled per-warp in issue_eligible_mask

    // Scheduler temporary variables (moved outside procedural block for synthesis)
    logic sched_found;
    int   sched_eligible_count;
    logic intra_hazard;

    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            rr_ptr <= 0;
            if_id[0].valid <= 0;
            if_id[1].valid <= 0;
            last_issued_valid <= 0;
            last_issued_warp <= 0;
            
            // Refactored State Reset
            for (int w=0; w<NUM_WARPS; w++) begin
                warp_pc[w]           <= 0;
                warp_state[w]        <= W_IDLE;
                warp_active_mask[w]  <= '1;
                warp_stack_ptr[w]    <= 0;
                warp_ret_ptr[w]      <= 0;
                warp_at_barrier[w] <= 0;
                warp_branch_tag[w]   <= 0;
            end
        end else begin
            // 1. Handle Branch Redirect (Highest Priority) - Independent of Stall
            if (cur_branch_taken) begin
                warp_pc[cur_branch_warp] <= cur_branch_target;
                // Flush Fetch Buffer if it matches flushed warp (even if stalled)
                if (if_id[0].valid && if_id[0].warp == cur_branch_warp) if_id[0].valid <= 0;
                if (if_id[1].valid && if_id[1].warp == cur_branch_warp) if_id[1].valid <= 0;
            end

            if (!stall_pipeline) begin
                if_id[0].valid <= 0;  // Default: Bubble
                if_id[1].valid <= 0;

                // 2. Kepler-Style Warp Selection (Select 1 warp, fetch PC and PC+1)
                if (!branch_taken_q && !cur_branch_taken) begin
                    logic warp_found;
                    logic [WARP_ID_WIDTH-1:0] selected_warp;
                    logic [63:0] inst_a, inst_b;
                    logic [7:0] pc_a, pc_b;
                    logic can_dual;
                    
                    warp_found = 0;
                    selected_warp = 0;
                    
                    // Round-robin search for eligible warp
                        
                    for (int i=0; i<NUM_WARPS; i++) begin
                        logic [WARP_ID_WIDTH-1:0] w;
                        w = (WARP_ID_WIDTH)'((32'(rr_ptr) + 32'(i)) % 32'(NUM_WARPS));
                        
                        if (issue_eligible_mask[w] && oc_dispatch_ready[0]) begin
                            selected_warp = w;
                            warp_found = 1;
                            break;
                        end else if (warp_state[w] == W_READY && cycle % 1000 == 0) begin
                             $display("CORE [%0t] SCHED_BLOCKED: Warp %0d Eligible=%b OC_Ready=%b", 
                                      $time, w, issue_eligible_mask[w], oc_dispatch_ready[0]);
                             scoreboard_diag(int'(w), prog_mem[w][ warp_pc[w][7:0] ]);
                        end
                    end
                    
                    if (warp_found) begin
                        pc_a = warp_pc[selected_warp][7:0];
                        pc_b = 8'(32'(pc_a) + 1);
                        
                        inst_a = prog_mem[selected_warp][pc_a];
                        inst_b = prog_mem[selected_warp][pc_b];
                        
                        // Always issue first instruction
                        if_id[0].valid <= 1;
                        if_id[0].warp  <= selected_warp;
                        if_id[0].pc    <= {24'b0, pc_a};
                        if_id[0].inst  <= inst_a;
                        if_id[0].branch_tag <= warp_branch_tag[selected_warp];
                        
                        // Check if we can dual-issue second instruction
                        // Intra-packet check: inst_b cannot depend on inst_a
                        begin : dual_hazard_check
                            opcode_t op_a, op_b;
                            logic [7:0] rd_a, rs1_b, rs2_b, rs3_b;
                            logic writes_a;
                            
                            op_a = opcode_t'(inst_a[63:56]);
                            op_b = opcode_t'(inst_b[63:56]);
                            rd_a = inst_a[55:48];
                            rs1_b = inst_b[47:40];
                            rs2_b = inst_b[39:32];
                            rs3_b = inst_b[27:20];
                            
                            // Check if inst_a writes to a register
                            writes_a = (op_a inside {OP_ADD,OP_SUB,OP_MUL,OP_IMAD,OP_SLT,OP_LDR,OP_MOV,OP_TID,
                                                   OP_FADD,OP_FSUB,OP_FMUL,OP_FDIV,OP_FFMA,OP_SFU_SIN,OP_SFU_COS,
                                                   OP_ITOF,OP_FTOI,OP_IDIV,OP_IREM,OP_AND,OP_OR,OP_XOR,OP_NOT,
                                                   OP_SHL,OP_SHR,OP_SHA,OP_ISETP,OP_FSETP,OP_LDS});
                            
                            intra_hazard = 0;
                            if (writes_a) begin
                                if (rd_a == rs1_b || rd_a == rs2_b || rd_a == rs3_b || rd_a == inst_b[55:48]) begin
                                    intra_hazard = 1;
                                end
                            end
                            
                            // Predicate RAW Hazard: inst_a writes Px, inst_b reads Px
                            if (op_a == OP_ISETP || op_a == OP_FSETP) begin
                                logic [2:0] pred_rd_a = inst_a[50:48];
                                if (inst_b[31:28] != 4'h7 && inst_b[30:28] == pred_rd_a) intra_hazard = 1; // Guard
                                if (op_b == OP_SELP && inst_b[2:0] == pred_rd_a) intra_hazard = 1;         // Source
                            end
                        end
                        
                        can_dual = can_dual_issue(inst_a, inst_b) && !intra_hazard && scoreboard_ok(int'(selected_warp), inst_b) && oc_dispatch_ready[1];
                        
                        if (can_dual) begin
                            // Dual-issue: Issue both instructions
                            if_id[1].valid <= 1;
                            if_id[1].warp  <= selected_warp;
                            if_id[1].pc    <= {24'b0, pc_b};
                            if_id[1].inst  <= inst_b;
                            if_id[1].branch_tag <= warp_branch_tag[selected_warp];
                            warp_pc[selected_warp] <= warp_pc[selected_warp] + 2;
                            
                            if (selected_warp == 0) begin
                                opcode_t op_a, op_b;
                                op_a = opcode_t'(inst_a[63:56]);
                                op_b = opcode_t'(inst_b[63:56]);
                                $display("CORE [%0t] KEPLER DUAL-ISSUE: Warp 0 PC=%h+%h Op=%s+%s", 
                                         $time, pc_a, pc_b, op_a.name(), op_b.name());
                            end
                        end else begin
                            // Single-issue: Only first instruction
                            if_id[1].valid <= 0;
                            warp_pc[selected_warp] <= warp_pc[selected_warp] + 1;
                            
                            if (selected_warp == 0) begin
                                opcode_t op_a;
                                op_a = opcode_t'(inst_a[63:56]);
                                $display("CORE [%0t] KEPLER SINGLE-ISSUE: Warp 0 PC=%h Op=%s", 
                                         $time, pc_a, op_a.name());
                            end
                        end
                        
                        // Update round-robin pointer
                        rr_ptr <= (32'(selected_warp) + 1) % 32'(NUM_WARPS);
                    end
                end
            end else begin
                 // STALL: Hold Pipeline State (Freeze IF/ID)
            end
        end
    end 
    //=========================================================================
    // PIPELINE STAGE: ID (Instruction Decode) - DUAL ISSUE
    //=========================================================================
    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            id_ex[0] <= '{op:OP_NOP, default:0};
            id_ex[1] <= '{op:OP_NOP, default:0};
            // Reset Scoreboard & Predicates here to be near reservation logic
            for (int w=0; w<NUM_WARPS; w++) begin
                warp_reg_writes[w] <= 0; 
                warp_pred_writes[w] <= 0; // Clear Predicate Scoreboard
                for (int l=0; l<WARP_SIZE; l++) preds[w][l] <= 0;
            end
            oc_wb_valid_q   <= 0;
            oc_wb_warp_q    <= 0;
            oc_wb_rd_q      <= 0;
            oc_wb_mask_q    <= 0;
            oc_wb_result_q  <= 0;
            oc_wb_we_q      <= 0;
            oc_wb_we_pred_q <= 0;
        end else begin
            // 1. Calculate Next State (Combinational Clear + Sequential Set)
            logic [NUM_REGS-1:0] next_sb [NUM_WARPS-1:0];
            logic [7:0]          next_pred_sb [NUM_WARPS-1:0];
            
            for (int w=0; w<NUM_WARPS; w++) begin
                // Start with current state, apply clears
                next_sb[w] = warp_reg_writes[w] & ~reg_clear_this_cycle[w];
                next_pred_sb[w] = warp_pred_writes[w] & ~pred_clear_this_cycle[w];
            end
            
            // Apply Predicate Updates (From Sync WB or Async MEM_RESP)
            if (oc_wb_valid[0] && oc_wb_we_pred_q[0]) begin
                 for (int l=0; l<WARP_SIZE; l++) begin
                     if (oc_wb_mask_q[0][l]) preds[oc_wb_warp_q[0]][l][oc_wb_rd_q[0][2:0]] <= oc_wb_result_q[0][l][0];
                 end
            end
            if (oc_wb_valid[1] && oc_wb_we_pred_q[1]) begin
                 for (int l=0; l<WARP_SIZE; l++) begin
                     if (oc_wb_mask_q[1][l]) preds[oc_wb_warp_q[1]][l][oc_wb_rd_q[1][2:0]] <= oc_wb_result_q[1][l][0];
                 end
            end

            // 2. Apply Sets if Pipeline Not Stalled
            if (!stall_pipeline) begin
                for (int p=0; p<2; p++) begin
                    if (if_id[p].valid) begin
                        opcode_t op;
                        op = opcode_t'(if_id[p].inst[63:56]);

                        // SECURITY: Do NOT set SB if instruction is Trash (Tag Mismatch)
                        if (if_id[p].branch_tag != warp_branch_tag[if_id[p].warp]) continue;
                        
                        // SECURITY: Do NOT set SB if instruction is currently being Flushed (Branch Taken NOW)
                        if (cur_branch_taken && cur_branch_warp == if_id[p].warp) continue;

                        if (op inside {OP_ADD,OP_SUB,OP_MUL,OP_IMAD,OP_SLT,OP_LDR,OP_MOV,OP_TID,
                                                           OP_FADD,OP_FSUB,OP_FMUL,OP_FDIV,OP_FTOI,
                                                           OP_SFU_SIN,OP_SFU_COS,OP_SFU_EX2,OP_SFU_LG2,
                                                           OP_SFU_RCP,OP_SFU_RSQ,OP_SFU_SQRT,OP_SFU_TANH,
                                                           OP_FFMA,
                                                           OP_IDIV,OP_IREM,
                                                           OP_IMIN,OP_IMAX,OP_IABS,
                                                           OP_FMIN,OP_FMAX,OP_FABS,
                                                           OP_AND,OP_OR,OP_XOR,OP_NOT,
                                                           OP_SHL,OP_SHR,OP_SHA,
                                                           OP_POPC,OP_CLZ,OP_BREV,OP_ITOF,
                                                           OP_NEG, OP_FNEG,
                                                           OP_CNOT,
                                                           OP_SLE,OP_SEQ,
                                                           OP_LDS}) begin
                            // Check for Branch Flush (Legacy Check - possibly redundant but safe)
                            if (!(branch_taken_q && branch_warp_q == if_id[p].warp)) begin
                                next_sb[if_id[p].warp][ 6'(if_id[p].inst[55:48]) ] = 1;
                            end
                        end
                        
                        // Set Predicate Scoreboard
                        if (op inside {OP_ISETP, OP_FSETP}) begin
                             if (!(branch_taken_q && branch_warp_q == if_id[p].warp)) begin
                                 next_pred_sb[if_id[p].warp][ if_id[p].inst[50:48] ] = 1; // RD is [2:0] for Pred Index
                             end
                        end
                    end
                end
                
                // Also handle other ID state updates (PC propagation etc)
                id_ex[0] <= '{op:OP_NOP, default:0};
                id_ex[1] <= '{op:OP_NOP, default:0};

                // Decode both instructions in parallel
                for (int p=0; p<2; p++) begin
                    if (if_id[p].valid) begin
                        opcode_t current_op;
                        current_op = opcode_t'(if_id[p].inst[63:56]);

                        // Check for Branch Flush (Shadow Instruction) or Tag Mismatch
                        if (if_id[p].branch_tag != warp_branch_tag[if_id[p].warp]) begin
                            // SQUASHED (Tag Mismatch)
                        end else begin
                            // Decode & Pass to OC
                            id_ex[p].valid <= 1;
                            id_ex[p].warp  <= if_id[p].warp;
                            id_ex[p].pc    <= if_id[p].pc;
                            id_ex[p].op    <= current_op;
                            id_ex[p].rd    <= if_id[p].inst[55:48];
                            id_ex[p].imm   <= {{12{if_id[p].inst[19]}}, if_id[p].inst[19:0]};
                            id_ex[p].pred_guard <= if_id[p].inst[31:28];
                            
                            // Read Source Predicate (ONLY For SELP) - With Bypass
                            if (current_op == OP_SELP) begin
                                for (int l=0; l<WARP_SIZE; l++) begin
                                     logic [2:0] p_idx;
                                     p_idx = if_id[p].inst[2:0];
                                     if (p_idx == 3'd7) begin
                                         id_ex[p].src_pred[l] <= 1'b1; // PT
                                     end else begin
                                         // Bypass from alu_wb (currently in WB stage)
                                         if (alu_wb.valid && alu_wb.we_pred && alu_wb.warp == if_id[p].warp && alu_wb.rd[2:0] == p_idx) begin
                                             id_ex[p].src_pred[l] <= alu_wb.result[l][0];
                                         end else begin
                                             id_ex[p].src_pred[l] <= preds[if_id[p].warp][l][p_idx]; 
                                         end
                                     end
                                end
                            end else begin
                                id_ex[p].src_pred <= '1; // Default to Always True for non-SELP ops
                            end
                            
                            id_ex[p].mask  <= warp_active_mask[if_id[p].warp];

                            // Pass register indices to OC
                            id_ex[p].rs1_idx <= if_id[p].inst[47:40];
                            id_ex[p].rs2_idx <= if_id[p].inst[39:32];
                            id_ex[p].rs3_idx <= if_id[p].inst[27:20];
                            
                            // Attach current Branch Tag
                            id_ex[p].branch_tag <= warp_branch_tag[if_id[p].warp];
                        end
                    end
                end
            end 
            
            // 3. Commit Scoreboard Update (Unconditionally)
            for (int w=0; w<NUM_WARPS; w++) begin
                warp_reg_writes[w] <= next_sb[w];
                warp_pred_writes[w] <= next_pred_sb[w];
            end
        end
    end

    // --- ID -> OC Dispatch wiring (Dual Issue) ---
    assign oc_dispatch_valid[0] = id_ex[0].valid;
    assign oc_dispatch_inst[0]  = id_ex[0];
    assign oc_dispatch_valid[1] = id_ex[1].valid;
    assign oc_dispatch_inst[1]  = id_ex[1];

    //=========================================================================
    // DISPATCH ROUTER: Route OC outputs to ALU or LSU Pipeline
    //=========================================================================
    // Instructions are routed to queues based on type (Memory vs Compute)
    // OC Ready signals (backpressure)
    // Prevent queues from growing infinitely. Stall OC if queues are full.
    // Use a conservative threshold (e.g., 8).
    // Signals for execution (Combinational from FIFO)
    id_ex_t alu_inst_exec;
    id_ex_t lsu_inst_exec;
    id_ex_t fpu_inst_exec;
    logic alu_valid_exec;
    logic lsu_valid_exec;
    logic fpu_valid_exec;
    
    // Internal FIFO Signals
    logic alu_push, lsu_push, fpu_push;
    logic alu_pop, lsu_pop, fpu_pop;
    id_ex_t alu_din, lsu_din, fpu_din;
    id_ex_t alu_dout, lsu_dout, fpu_dout; 
    logic alu_full, lsu_full, fpu_full;
    logic alu_empty, lsu_empty, fpu_empty;
    int alu_count, lsu_count, fpu_count;

    // ------------------------------------------------------------------------
    // INSTANTIATE FIFOs (DEPTH 8)
    // ------------------------------------------------------------------------
    fifo #( .DEPTH(8), .T(id_ex_t) ) alu_fifo (
        .clk(clk), .rst_n(rst_n),
        .push(alu_push), .pop(alu_pop),
        .data_in(alu_din),
        .data_out(alu_dout), // Combinational Peek
        .full(alu_full), .empty(alu_empty), .count(alu_count)
    );

    fifo #( .DEPTH(8), .T(id_ex_t) ) lsu_fifo (
        .clk(clk), .rst_n(rst_n),
        .push(lsu_push), .pop(lsu_pop),
        .data_in(lsu_din),
        .data_out(lsu_dout), 
        .full(lsu_full), .empty(lsu_empty), .count(lsu_count)
    );

    fifo #( .DEPTH(8), .T(id_ex_t) ) fpu_fifo (
        .clk(clk), .rst_n(rst_n),
        .push(fpu_push), .pop(fpu_pop),
        .data_in(fpu_din),
        .data_out(fpu_dout), 
        .full(fpu_full), .empty(fpu_empty), .count(fpu_count)
    );

    // ------------------------------------------------------------------------
    // CONSUMER LOGIC (Combinational Ready/Valid/Pop)
    // ------------------------------------------------------------------------
    // Validate Execution Input: Valid ONLY if FIFO has data
    assign alu_valid_exec = !alu_empty;
    // LSU Gating: Never launch if no TX ID is available (prevents $fatal in MEM)
    assign lsu_valid_exec = !lsu_empty && 
                           !((lsu_dout.op == OP_LDR || lsu_dout.op == OP_STR || lsu_dout.op == OP_LDS || lsu_dout.op == OP_STS) && 
                             tx_id_fifo_empty[lsu_dout.warp]);
    assign fpu_valid_exec = !fpu_empty;
    
    // Assign Execution Instruction: Directly from FIFO peek (or NOP if empty)
    assign alu_inst_exec = alu_valid_exec ? alu_dout : '{op:OP_NOP, default:0};
    assign lsu_inst_exec = lsu_valid_exec ? lsu_dout : '{op:OP_NOP, default:0};
    assign fpu_inst_exec = fpu_valid_exec ? fpu_dout : '{op:OP_NOP, default:0};

    // Auto-Pop Logic: Pop from FIFOs when valid
    logic alu_can_commit;
    assign alu_pop = alu_valid_exec && alu_can_commit;
    
    // LSU Pop logic: Only advance if the MEM stage can accept a new instruction
    logic lsu_mem_consumed;
    assign lsu_pop = lsu_valid_exec && (!lsu_mem.valid || lsu_mem_consumed);

    // FPU Pop logic with explicit backpressure from Writeback Arbiter
    logic stall_fpu_wb;
    assign fpu_pop = fpu_valid_exec && !stall_pipeline && !stall_fpu_wb;

    // ------------------------------------------------------------------------
    // PRODUCER LOGIC (Push to FIFOs)
    // ------------------------------------------------------------------------
    // Router logic: Determine which FIFO to push instructions based on unit type
    
    always_comb begin
        alu_push = 0;
        lsu_push = 0;
        fpu_push = 0;
        alu_din = '{op:OP_NOP, default:0};
        lsu_din = '{op:OP_NOP, default:0};
        fpu_din = '{op:OP_NOP, default:0};
        oc_ex_ready = 2'b00;
        
        // 1. Check Port 0
        if (oc_ex_valid[0]) begin
            case (get_unit_type(oc_ex_inst[0].op))
                UNIT_LSU: begin
                    if (!lsu_full || lsu_pop) begin
                        lsu_push = 1; lsu_din = oc_ex_inst[0];
                        oc_ex_ready[0] = 1;
                        // $display("CORE [%0t] ROUTER_P0: LSU Push Op=%s", $time, oc_ex_inst[0].op.name());
                    end
                end
                UNIT_FPU: begin
                     if (!fpu_full || fpu_pop) begin
                        fpu_push = 1; fpu_din = oc_ex_inst[0];
                        oc_ex_ready[0] = 1;
                    end
                end
                default: begin // ALU, CTRL
                     // ALU is coupled to stall_pipeline, so we cannot use prediction here (creates loop)
                     if (!alu_full) begin
                        alu_push = 1; alu_din = oc_ex_inst[0];
                        oc_ex_ready[0] = 1;
                        $display("CORE [%0t] ROUTER_P0: ALU Push Warp=%0d PC=%h Op=%s", $time, oc_ex_inst[0].warp, oc_ex_inst[0].pc, oc_ex_inst[0].op.name());
                    end
                end
            endcase
        end
        
        // 2. Check Port 1 (Prioritize if FIFO available)
        if (oc_ex_valid[1]) begin
             case (get_unit_type(oc_ex_inst[1].op))
                UNIT_LSU: begin
                    if (!lsu_push && (!lsu_full || lsu_pop)) begin
                        lsu_push = 1; lsu_din = oc_ex_inst[1];
                        oc_ex_ready[1] = 1;
                    end
                end
                UNIT_FPU: begin
                     if (!fpu_push && (!fpu_full || fpu_pop)) begin
                        fpu_push = 1; fpu_din = oc_ex_inst[1];
                        oc_ex_ready[1] = 1;
                    end
                end
                default: begin // ALU
                     if (!alu_push && !alu_full) begin
                        alu_push = 1; alu_din = oc_ex_inst[1];
                        oc_ex_ready[1] = 1;
                        $display("CORE [%0t] ROUTER_P1: ALU Push Warp=%0d PC=%h Op=%s", $time, oc_ex_inst[1].warp, oc_ex_inst[1].pc, oc_ex_inst[1].op.name());
                    end
                end
            endcase
        end

        // ASSERTION: The dual-issue scheduler (can_dual_issue) must prevent structural hazards.
        // If we reach here and both ports target the same backend resource, it is a design bug.
    end

    // Logging (Moved to separate always_ff to avoid clutter in comb block)
    always_ff @(posedge clk) begin
       if (alu_push && alu_din.warp == 0) 
            $display("CORE [%0t] ROUTER: Warp 0 Op=%s -> ALU FIFO (Combinational Push)", $time, alu_din.op.name());
       if (lsu_push && lsu_din.warp == 0) 
            $display("CORE [%0t] ROUTER: Warp 0 Op=%s -> LSU FIFO (Combinational Push)", $time, lsu_din.op.name());
       
       // Debug to catch Phantom LSU Pushes
       if (oc_ex_valid[0] && oc_ex_inst[0].warp == 0 && !alu_push && !lsu_push && !fpu_push)
            $display("CORE [%0t] ROUTER: Warp 0 Dropped? Op=%s Unit=%0d", $time, oc_ex_inst[0].op.name(), get_unit_type(oc_ex_inst[0].op));
       if (lsu_push && get_unit_type(lsu_din.op) != UNIT_LSU)
            $display("CORE [%0t] ROUTER ERROR: Pushing Non-LSU Op %s to LSU FIFO!", $time, lsu_din.op.name());
       if (!lsu_empty && !lsu_pop && !lsu_push)
            $display("CORE [%0t] LSU FIFO STATE: Count=%0d HeadOp=%s", $time, lsu_count, lsu_dout.op.name());
    end

    //=========================================================================
    // PIPELINE STAGE: EX (Execute)
    //=========================================================================
    // - Performs ALU operations (ADD, SUB, MUL, SLT)
    // - Resolves branches and updates divergence stack
    // - Calculates memory addresses for loads/stores
    // - Handles thread divergence (BEQ/BNE) and reconvergence (JOIN)
    //=========================================================================
    
    // ------------------------------------------------------------------------
    // Execution Mask Logic (Combinational) - Handles Predication & Forwarding
    // ------------------------------------------------------------------------
    logic [WARP_SIZE-1:0] exec_mask_alu;
    logic [WARP_SIZE-1:0] exec_mask_lsu;
    logic [WARP_SIZE-1:0] exec_mask_fpu;
    
    // ALU Execution Mask
    always_comb begin
        logic [WARP_SIZE-1:0] p_vals;
        logic [2:0] p_id;
        logic p_neg;
        
        exec_mask_alu = 0;
        
        if (alu_valid_exec) begin
            p_id = alu_inst_exec.pred_guard[2:0];
            p_neg = alu_inst_exec.pred_guard[3];

            for (int l=0; l<WARP_SIZE; l++) begin
                p_vals[l] = 0;
                if (p_id == 7) begin
                    p_vals[l] = 1'b1; // PT (Always True)
                end else begin
                    // Forwarding from ALU WB (Current WB stage)
                    if (alu_wb.valid && alu_wb.we_pred && alu_wb.warp == alu_inst_exec.warp && alu_wb.rd[2:0] == p_id) begin
                         p_vals[l] = alu_wb.result[l][0];
                    end 
                    // Forwarding from Async MEM WB
                    else if (mem_resp_wb.valid && mem_resp_wb.we_pred && mem_resp_wb.warp == alu_inst_exec.warp && mem_resp_wb.rd[2:0] == p_id) begin
                         p_vals[l] = mem_resp_wb.result[l][0];
                    end else begin
                         p_vals[l] = preds[alu_inst_exec.warp][l][p_id];
                    end
                end
                // CRITICAL: Use current architectural active_mask to handle divergence correctly
                exec_mask_alu[l] = alu_inst_exec.mask[l] & (p_neg ? ~p_vals[l] : p_vals[l]);
            end
        end
    end
    
    // LSU Execution Mask
    always_comb begin
        logic [WARP_SIZE-1:0] p_vals;
        logic [2:0] p_id;
        logic p_neg;
        
        exec_mask_lsu = 0;
        
        if (lsu_valid_exec) begin
            p_id = lsu_inst_exec.pred_guard[2:0];
            p_neg = lsu_inst_exec.pred_guard[3];

            for (int l=0; l<WARP_SIZE; l++) begin
                p_vals[l] = 0;
                if (p_id == 7) begin
                    p_vals[l] = 1'b1; 
                end else begin
                    if (alu_wb.valid && alu_wb.we_pred && alu_wb.warp == lsu_inst_exec.warp && alu_wb.rd[2:0] == p_id) begin
                         p_vals[l] = alu_wb.result[l][0];
                    end else if (mem_resp_wb.valid && mem_resp_wb.we_pred && mem_resp_wb.warp == lsu_inst_exec.warp && mem_resp_wb.rd[2:0] == p_id) begin
                         p_vals[l] = mem_resp_wb.result[l][0];
                    end else begin
                         p_vals[l] = preds[lsu_inst_exec.warp][l][p_id];
                    end
                end
                // CRITICAL: Use the mask dispatched with the instruction
                exec_mask_lsu[l] = lsu_inst_exec.mask[l] & (p_neg ? ~p_vals[l] : p_vals[l]);
            end
        end
    end
    
    // Branch evaluation moved to EX stage sequential block

    // FPU Execution Mask
    always_comb begin
        logic [WARP_SIZE-1:0] p_vals;
        logic [2:0] p_id;
        logic p_neg;
        
        exec_mask_fpu = 0;
        
        if (fpu_valid_exec) begin
            p_id = fpu_inst_exec.pred_guard[2:0];
            p_neg = fpu_inst_exec.pred_guard[3];

            for (int l=0; l<WARP_SIZE; l++) begin
                p_vals[l] = 0;
                if (p_id == 7) begin
                    p_vals[l] = 1'b1; 
                end else begin
                    if (alu_wb.valid && alu_wb.we_pred && alu_wb.warp == fpu_inst_exec.warp && alu_wb.rd[2:0] == p_id) begin
                         p_vals[l] = alu_wb.result[l][0];
                    end else if (mem_resp_wb.valid && mem_resp_wb.we_pred && mem_resp_wb.warp == fpu_inst_exec.warp && mem_resp_wb.rd[2:0] == p_id) begin
                         p_vals[l] = mem_resp_wb.result[l][0];
                    end else begin
                         p_vals[l] = preds[fpu_inst_exec.warp][l][p_id];
                    end
                end
                // CRITICAL: Use the mask dispatched with the instruction
                exec_mask_fpu[l] = fpu_inst_exec.mask[l] & (p_neg ? ~p_vals[l] : p_vals[l]);
            end
        end
    end

    // ------------------------------------------------------------------------
    // FPU Instantiation (32 Lanes)
    // ------------------------------------------------------------------------
    logic [WARP_SIZE-1:0][31:0] fpu_out;
    logic [3:0] fpu_op_code;
    
    // Simple Opcode Decoder for FPU
    always_comb begin
        case (fpu_inst_exec.op)
            OP_FADD: fpu_op_code = 4'd10; // Add
            OP_FSUB: fpu_op_code = 4'd3;  // Sub
            OP_FMUL: fpu_op_code = 4'd1;  // Mul
            OP_FDIV: fpu_op_code = 4'd2;  // Div
            OP_FTOI: fpu_op_code = 4'd9;  // Float -> Int
            OP_ITOF: fpu_op_code = 4'd12; // Int -> Float
            default: fpu_op_code = 4'd10;
        endcase
    end

    // Lane Generation for FPU
    genvar k;
    generate
        for (k=0; k<WARP_SIZE; k++) begin : fpu_lane
            // Wires for exceptions (ignored for now)
            wire fpu_exc, fpu_ovf, fpu_unf;
            
            ALU fpu_inst (
                .a_operand(fpu_en ? fpu_inst_exec.rs1[k] : 32'b0),
                .b_operand(fpu_en ? fpu_inst_exec.rs2[k] : 32'b0),
                .Operation(fpu_op_code),
                .ALU_Output(fpu_out[k]),
                .Exception(fpu_exc),
                .Overflow(fpu_ovf),
                .Underflow(fpu_unf)
            );
        end
    endgenerate

    // ------------------------------------------------------------------------
    // SFU Instantiation (32 Lanes)
    // ------------------------------------------------------------------------
    logic [WARP_SIZE-1:0][15:0] sfu_out;
    sfu_op_t sfu_op_code;

    // SFU Operation Decoder
    always_comb begin
        case (fpu_inst_exec.op)
            OP_SFU_SIN:  sfu_op_code = SFU_SIN;
            OP_SFU_COS:  sfu_op_code = SFU_COS;
            OP_SFU_EX2:  sfu_op_code = SFU_EX2;
            OP_SFU_LG2:  sfu_op_code = SFU_LG2;
            OP_SFU_RCP:  sfu_op_code = SFU_RCP;
            OP_SFU_RSQ:  sfu_op_code = SFU_RSQ;
            OP_SFU_SQRT: sfu_op_code = SFU_SQRT;
            OP_SFU_TANH: sfu_op_code = SFU_TANH;
            default:     sfu_op_code = SFU_SIN; 
        endcase
    end

    // Lane Generation for SFU
    genvar m;
    generate
        for (m=0; m<WARP_SIZE; m++) begin : sfu_lane
            sfu_single_cycle #(.LUT_SIZE(256)) sfu_inst (
                .operation(sfu_op_code),
                .operand(sfu_en ? fpu_inst_exec.rs1[m][15:0] : 16'b0), // Gated
                .result(sfu_out[m])
            );
        end
    endgenerate

    // Lane Generation for FMA
    logic [WARP_SIZE-1:0][31:0] fma_out;
    logic [WARP_SIZE-1:0] fma_exception; // Unused for now
    
    // Mutual Exclusion Enables
    logic fpu_en, sfu_en, fma_en;
    always_comb begin
        fpu_en = 0; sfu_en = 0; fma_en = 0;
        if (fpu_valid_exec) begin
            if (fpu_inst_exec.op >= OP_SFU_SIN && fpu_inst_exec.op <= OP_SFU_TANH) sfu_en = 1;
            else if (fpu_inst_exec.op == OP_FFMA || fpu_inst_exec.op == OP_FADD || fpu_inst_exec.op == OP_FMUL) fma_en = 1;
            else fpu_en = 1;
        end
    end

    // Helper signals for FMA operands
    logic [WARP_SIZE-1:0][31:0] fma_op_a;
    logic [WARP_SIZE-1:0][31:0] fma_op_b;
    logic [WARP_SIZE-1:0][31:0] fma_op_c;

    always_comb begin 
        for(int i=0; i<WARP_SIZE; i++) begin
            // Default: FFMA (A * B + C)
            fma_op_a[i] = fpu_inst_exec.rs1[i];
            fma_op_b[i] = fpu_inst_exec.rs2[i];
            fma_op_c[i] = fpu_inst_exec.rs3[i]; 

            // Special cases
            if (fpu_inst_exec.op == OP_FADD) begin
                // A + B -> Use (A * 1.0) + B
                fma_op_a[i] = fpu_inst_exec.rs1[i];
                fma_op_b[i] = 32'h3F800000; // 1.0
                fma_op_c[i] = fpu_inst_exec.rs2[i]; 
            end else if (fpu_inst_exec.op == OP_FMUL) begin
                // A * B -> Use (A * B) + 0.0
                fma_op_a[i] = fpu_inst_exec.rs1[i];
                fma_op_b[i] = fpu_inst_exec.rs2[i]; 
                fma_op_c[i] = 32'h00000000; // 0.0
            end 
            // Actually usually handled by negating operand B logic or separate Sub unit.
            // For now let's just fix FADD/FMUL.
        end 
    end

    genvar f;
    generate
        for (f=0; f<WARP_SIZE; f++) begin : fma_lane
            FMA fma_inst (
                .a_operand(fma_en ? fma_op_a[f] : 32'b0),
                .b_operand(fma_en ? fma_op_b[f] : 32'b0),
                .c_operand(fma_en ? fma_op_c[f] : 32'b0),
                .result(fma_out[f]),
                .Exception(fma_exception[f])
            );
        end
    endgenerate

    // 2. Separate Execution Paths (ALU/Compute vs LSU/Memory)
    
    // ------------------------------------------------------------------------
    // Integer ALU Instantiation (Combinational)
    // ------------------------------------------------------------------------
    logic [WARP_SIZE-1:0][31:0] int_alu_out;
    logic [WARP_SIZE-1:0][31:0] sfu_out_32b;
    
    // Sign-extend SFU output to 32 bits (fixed point 1.15)
    generate 
        for(genvar i=0; i<WARP_SIZE; i++) assign sfu_out_32b[i] = {{16{sfu_out[i][15]}}, sfu_out[i]};
    endgenerate

    // Re-calculate src_pred in EX stage for SELP bypass
    logic [WARP_SIZE-1:0] alu_inst_exec_src_pred;
    always_comb begin
        for (int l=0; l<WARP_SIZE; l++) begin
            logic [2:0] p_idx;
            p_idx = alu_inst_exec.imm[2:0]; // PredID for SELP is in imm[2:0]
            if (p_idx == 7) begin
                alu_inst_exec_src_pred[l] = 1'b1;
            end else begin
                if (alu_wb.valid && alu_wb.we_pred && alu_wb.warp == alu_inst_exec.warp && alu_wb.rd[2:0] == p_idx) begin
                    alu_inst_exec_src_pred[l] = alu_wb.result[l][0];
                end else if (mem_resp_wb.valid && mem_resp_wb.we_pred && mem_resp_wb.warp == alu_inst_exec.warp && mem_resp_wb.rd[2:0] == p_idx) begin
                    alu_inst_exec_src_pred[l] = mem_resp_wb.result[l][0];
                end else begin
                    alu_inst_exec_src_pred[l] = preds[alu_inst_exec.warp][l][p_idx];
                end
            end
        end
    end

    int_alu i_alu_inst (
        .op(alu_inst_exec.op),
        .imm(alu_inst_exec.imm),
        .rs1(alu_inst_exec.rs1),
        .rs2(alu_inst_exec.rs2),
        .rs3(alu_inst_exec.rs3),
        .src_pred(alu_inst_exec.op == OP_SELP ? alu_inst_exec_src_pred : alu_inst_exec.src_pred),
        
        .warp(alu_inst_exec.warp),
        .result(int_alu_out)
    );
    
    // ------------------------------------------------------------------------
    // PATH A: ALU / Compute Pipeline (Single Cycle Execution)
    // ------------------------------------------------------------------------
    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            alu_wb <= '{op:OP_NOP, valid:0, src:WB_ALU, warp:0, rd:0, mask:0, result:0, we:0, we_pred:0};
        end else begin
            alu_wb <= '{op:OP_NOP, valid:0, src:WB_ALU, warp:0, rd:0, mask:0, result:0, we:0, we_pred:0};
            
            if (alu_valid_exec) begin
                // Process ALU instruction
                $display("CORE [%0t] ALU EXEC: Warp=%0d PC=%h Op=%s Mask=%h Res0=%h Res16=%h", 
                    $time, alu_inst_exec.warp, alu_inst_exec.pc, alu_inst_exec.op.name(), exec_mask_alu, int_alu_out[0], int_alu_out[16]);
                
                // Check for Branch Flush (Tag Mismatch)
                if (alu_inst_exec.branch_tag != warp_branch_tag[alu_inst_exec.warp]) begin
                    // SQUASHED: We must still progress to WB to clear scoreboard entry for 'rd'
                    alu_wb.valid <= 1;
                    alu_wb.src   <= WB_ALU;
                    alu_wb.warp  <= alu_inst_exec.warp;
                    alu_wb.op    <= OP_NOP;
                    alu_wb.rd    <= alu_inst_exec.rd;
                    alu_wb.mask  <= 0;
                    alu_wb.we    <= 0;
                    alu_wb.we_pred <= 0;
                    alu_wb.result <= 0;
                end else if (branch_taken_q && branch_warp_q == alu_inst_exec.warp) begin
                    // Legacy flush (Shadow instruction case)
                    alu_wb.valid <= 1;
                    alu_wb.src   <= WB_ALU;
                    alu_wb.warp  <= alu_inst_exec.warp;
                    alu_wb.op    <= OP_NOP;
                    alu_wb.rd    <= alu_inst_exec.rd;
                    alu_wb.mask  <= 0;
                    alu_wb.we    <= 0;
                    alu_wb.we_pred <= 0;
                    alu_wb.result <= 0;
                end else begin
                    // Valid Execution
                    alu_wb.valid <= 1;
                    alu_wb.src   <= WB_ALU;
                    alu_wb.warp  <= alu_inst_exec.warp;
                    alu_wb.op    <= alu_inst_exec.op;
                    alu_wb.rd    <= alu_inst_exec.rd;
                    alu_wb.mask  <= exec_mask_alu;
                    
                    // Set Write Enable for standard compute ops
                    if (alu_inst_exec.op != OP_BRA && alu_inst_exec.op != OP_BEQ && 
                        alu_inst_exec.op != OP_BNE && alu_inst_exec.op != OP_EXIT &&
                        alu_inst_exec.op != OP_BAR && alu_inst_exec.op != OP_SSY &&
                        alu_inst_exec.op != OP_JOIN) begin
                        alu_wb.we <= 1;
                    end else begin
                        alu_wb.we <= 0;
                    end

                    // Set Predicate Write Enable
                    if (alu_inst_exec.op == OP_ISETP || alu_inst_exec.op == OP_FSETP) begin
                        alu_wb.we_pred <= 1;
                    end else begin
                        alu_wb.we_pred <= 0;
                    end
                    
                    
                    // Unified Result Writeback (from int_alu)
                    alu_wb.result <= int_alu_out;

                    // Control Flow Side-Effects (State Updates)
                    case (alu_inst_exec.op)
                        OP_SSY: begin
                            if (|exec_mask_alu) begin
                                stack_pc[alu_inst_exec.warp][ 5'(warp_stack_ptr[alu_inst_exec.warp]) ]   <= alu_inst_exec.pc + alu_inst_exec.imm;
                                stack_mask[alu_inst_exec.warp][ 5'(warp_stack_ptr[alu_inst_exec.warp]) ] <= warp_active_mask[alu_inst_exec.warp];
                                warp_stack_ptr[alu_inst_exec.warp] <= warp_stack_ptr[alu_inst_exec.warp] + 1;
                                $display("STACK [%0t] PUSH: Warp %0d Ptr %0d PC %h Mask %h", $time, alu_inst_exec.warp, warp_stack_ptr[alu_inst_exec.warp], alu_inst_exec.pc + alu_inst_exec.imm, warp_active_mask[alu_inst_exec.warp]);
                            end
                        end
                        OP_JOIN: begin
                            if (warp_stack_ptr[alu_inst_exec.warp] > 0) begin
                                warp_active_mask[alu_inst_exec.warp] <= stack_mask[alu_inst_exec.warp][ 5'(warp_stack_ptr[alu_inst_exec.warp] - 1) ];
                                warp_stack_ptr[alu_inst_exec.warp] <= warp_stack_ptr[alu_inst_exec.warp] - 1;
                            end
                        end
                        OP_BAR: begin
                            if (!barrier_active) begin
                                barrier_expected <= '0;
                                for (int i = 0; i < NUM_WARPS; i++) begin
                                    if (warp_state[i] == W_READY || warp_state[i] == W_BARRIER) barrier_expected[i] <= 1;
                                end
                                barrier_active <= 1;
                                barrier_initialized <= 0;
                            end
                            if (barrier_seen_epoch[alu_inst_exec.warp] != barrier_epoch) begin
                                barrier_seen_epoch[alu_inst_exec.warp] <= barrier_epoch;
                                barrier_mask[alu_inst_exec.warp]       <= 1'b1;
                            end
                            if (barrier_active && !barrier_initialized) barrier_initialized <= 1;
                            if (barrier_initialized && 
                                ((barrier_mask | (1 << alu_inst_exec.warp)) & barrier_expected) == barrier_expected && barrier_expected != 0) begin
                                barrier_mask        <= '0;
                                barrier_epoch       <= ~barrier_epoch;
                                barrier_seen_epoch  <= '0;
                                barrier_active      <= 0;
                                barrier_initialized <= 0;
                            end
                        end
                        OP_CALL: begin
                            ret_stack[alu_inst_exec.warp][ 3'(warp_ret_ptr[alu_inst_exec.warp]) ] <= alu_inst_exec.pc + 1;
                            warp_ret_ptr[alu_inst_exec.warp] <= warp_ret_ptr[alu_inst_exec.warp] + 1;
                        end
                        OP_RET: begin
                            if (warp_ret_ptr[alu_inst_exec.warp] > 0) begin
                                warp_ret_ptr[alu_inst_exec.warp] <= warp_ret_ptr[alu_inst_exec.warp] - 1;
                            end
                        end
                        OP_BEQ, OP_BNE: begin
                            logic [WARP_SIZE-1:0] taken_mask;
                            logic any_taken, any_not_taken;
                            taken_mask = 0;
                            for (int l=0; l<WARP_SIZE; l++) begin
                                if (exec_mask_alu[l]) begin
                                     logic eq;
                                     eq = (alu_inst_exec.rs1[l] == alu_inst_exec.rs2[l]);
                                     if ((alu_inst_exec.op == OP_BEQ && eq) || (alu_inst_exec.op == OP_BNE && !eq)) taken_mask[l] = 1;
                                end
                            end
                            any_taken = |taken_mask;
                            any_not_taken = |(exec_mask_alu & ~taken_mask);
                            if (alu_inst_exec.warp == 0) begin
                                $display("CORE [%0t] BEQ: PC=%h Mask=%h Taken=%h AnyT=%b AnyNT=%b", 
                                    $time, alu_inst_exec.pc, exec_mask_alu, taken_mask, any_taken, any_not_taken);
                            end
                            if (any_taken && any_not_taken) begin
                                // Divergence Side-Effect
                                stack_pc[alu_inst_exec.warp][ 5'(warp_stack_ptr[alu_inst_exec.warp]) ] <= alu_inst_exec.pc + 1;
                                stack_mask[alu_inst_exec.warp][ 5'(warp_stack_ptr[alu_inst_exec.warp]) ] <= (exec_mask_alu & ~taken_mask);
                                warp_stack_ptr[alu_inst_exec.warp] <= warp_stack_ptr[alu_inst_exec.warp] + 1;
                                warp_active_mask[alu_inst_exec.warp] <= taken_mask;
                            end
                        end
                        default: ;
                    endcase
                end
            end
            
            // Update Tag on Branch Taken
            if (cur_branch_taken && alu_can_commit) begin
                warp_branch_tag[cur_branch_warp] <= warp_branch_tag[cur_branch_warp] + 1;
            end
        end
    end

    // ALU Commit Logic: Define when an executed instruction can actually retire
    always_comb begin
        alu_can_commit = 1;
        if (alu_valid_exec && (alu_inst_exec.branch_tag == warp_branch_tag[alu_inst_exec.warp])) begin
            case (alu_inst_exec.op)
                OP_BAR, OP_EXIT: begin
                    int w = int'(alu_inst_exec.warp);
                    logic lsu_pipeline_busy;
                    lsu_pipeline_busy = (mshr_count[w] != 0) || 
                                       (lsu_valid_exec && lsu_inst_exec.warp == alu_inst_exec.warp) ||
                                       (lsu_mem.valid && lsu_mem.warp == alu_inst_exec.warp);
                    if (lsu_pipeline_busy)
                        alu_can_commit = 0;
                end
                default: alu_can_commit = 1;
            endcase
        end
    end

    // COMBINATIONAL BRANCH DETERMINATION
    always_comb begin
        cur_branch_taken  = 0;
        cur_branch_target = 0;
        cur_branch_warp   = 0;

        if (alu_valid_exec && (alu_inst_exec.branch_tag == warp_branch_tag[alu_inst_exec.warp])) begin
            case (alu_inst_exec.op)
                OP_BRA: begin
                    if (|exec_mask_alu) begin
                        cur_branch_taken = 1;
                        cur_branch_target = alu_inst_exec.pc + alu_inst_exec.imm;
                        cur_branch_warp = alu_inst_exec.warp;
                    end
                end
                OP_BEQ, OP_BNE: begin
                    if (|exec_mask_alu) begin
                        logic [WARP_SIZE-1:0] taken_mask;
                        for (int l=0; l<WARP_SIZE; l++) begin
                            logic eq;
                            eq = (alu_inst_exec.rs1[l] == alu_inst_exec.rs2[l]);
                            taken_mask[l] = (alu_inst_exec.op == OP_BEQ ? eq : !eq);
                        end
                        if (| (exec_mask_alu & taken_mask)) begin
                            cur_branch_taken = 1;
                            cur_branch_target = alu_inst_exec.pc + alu_inst_exec.imm;
                            cur_branch_warp = alu_inst_exec.warp;
                        end
                    end
                end
                OP_CALL: begin
                    cur_branch_taken = 1;
                    cur_branch_target = alu_inst_exec.pc + alu_inst_exec.imm;
                    cur_branch_warp = alu_inst_exec.warp;
                end
                OP_RET: begin
                    if (warp_ret_ptr[alu_inst_exec.warp] > 0) begin
                        cur_branch_taken = 1;
                        cur_branch_target = ret_stack[alu_inst_exec.warp][ 3'(warp_ret_ptr[alu_inst_exec.warp] - 1) ];
                        cur_branch_warp = alu_inst_exec.warp;
                    end
                end
                OP_EXIT: begin
                    cur_branch_taken = 1;
                    cur_branch_target = alu_inst_exec.pc;
                    cur_branch_warp = alu_inst_exec.warp;
                end
                OP_JOIN: begin
                    if (warp_stack_ptr[alu_inst_exec.warp] > 0) begin
                        cur_branch_taken  = 1;
                        cur_branch_target = stack_pc[alu_inst_exec.warp][ 5'(warp_stack_ptr[alu_inst_exec.warp] - 1) ];
                        cur_branch_warp   = alu_inst_exec.warp;
                    end
                end
                OP_SSY: begin
                    if (|exec_mask_alu) begin
                        cur_branch_taken  = 1;
                        cur_branch_target = alu_inst_exec.pc + 1;
                        cur_branch_warp   = alu_inst_exec.warp;
                    end
                end
                default: ;
            endcase
        end
    end

    // ------------------------------------------------------------------------
    // PATH B: LSU / Memory Pipeline (Address Calculation)
    // ------------------------------------------------------------------------
    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            lsu_mem <= '{op:OP_NOP, valid:0, warp:0, rd:0, mask:0, addresses:0, store_data:0, default:0};
        end else begin
            if (lsu_mem_consumed || !lsu_mem.valid) begin
                // Load Next from FIFO or clear
                lsu_mem <= '{op:OP_NOP, valid:0, warp:0, rd:0, mask:0, addresses:0, store_data:0, default:0};
                
                if (lsu_valid_exec) begin
                    if (lsu_inst_exec.branch_tag != warp_branch_tag[lsu_inst_exec.warp]) begin 
                        // SQUASHED: Emit "Shadow NOP" to clear scoreboard in WB stage
                        lsu_mem <= '{
                            op: OP_NOP,
                            valid: 1,      // KEEP VALID so it flows to WB
                            warp: lsu_inst_exec.warp,
                            rd: lsu_inst_exec.rd, // Preserve RD for scoreboard clear
                            mask: '0,      // Mask 0 = No Side Effects
                            addresses: 0,
                            store_data: 0,
                            default: 0
                        }; 
                    end else begin
                        // Valid Execution
                        lsu_mem.valid <= 1;
                        lsu_mem.warp  <= lsu_inst_exec.warp;
                        lsu_mem.op    <= lsu_inst_exec.op;
                        lsu_mem.rd    <= lsu_inst_exec.rd;
                        lsu_mem.mask  <= exec_mask_lsu;
                        
                        // Address Calculation (LDR/STR)
                        for (int l=0; l<WARP_SIZE; l++) begin
                            lsu_mem.addresses[l] <= lsu_inst_exec.rs1[l] + lsu_inst_exec.imm;
                            lsu_mem.store_data[l] <= lsu_inst_exec.rs2[l];
                        end
                    end
                end
            end
        end
    end
    
    // ------------------------------------------------------------------------
    // PIPELINE STAGE: MEM (Memory Access)
    // ------------------------------------------------------------------------
    // - Issues load/store requests to L1 cache (non-blocking)
    // - Allocates transaction IDs from free pool for tracking
    // - Stores request metadata in MSHR table for async completion
    // - Coalesces memory accesses across threads in a warp
    //=========================================================================
    
    // Signals for Memory Subsystem
    logic mem_busy;
    logic coalescer_valid;
    logic l1_req_valid, l1_req_rw, l1_req_ready, l1_resp_valid;
    logic [31:0] l1_req_addr;
    logic [1023:0] l1_req_wdata;
    logic [1023:0] l1_resp_rdata; // Defined as logic
    logic [WARP_SIZE-1:0] l1_req_mask;

    // ========================================================================
    // LSU REPLAY MECHANISM (Uncoalesced Access Handling)
    // ========================================================================
    
    // Replay Queue Entry Structure
    typedef struct packed {
        logic valid;
        logic [WARP_SIZE-1:0] pending_mask;
        logic [7:0] warp;
        logic [7:0] rd;
        logic [7:0] op;
        logic [WARP_SIZE-1:0][31:0] addresses;
        logic [WARP_SIZE-1:0][31:0] store_data;
    } replay_entry_t;
    
    // Per-warp replay queue (one entry per warp)
    replay_entry_t replay_queue [NUM_WARPS];
    
    // Replay arbiter signals
    logic [NUM_WARPS-1:0] replay_valid;
    logic [WARP_ID_WIDTH-1:0] replay_granted_warp;
    logic replay_grant_valid;
    
    // Current request source (new LSU or replay)
    lsu_mem_t current_lsu_request;
    logic current_is_replay;
    
    // Split calculation signals
    logic [WARP_SIZE-1:0] current_split_mask;
    logic [WARP_SIZE-1:0] next_split_mask;
    logic split_is_last;
    int   split_leader;
    logic mem_request_valid;
    
    // Helper to find first active lane
    function automatic int get_first_active_lane(logic [WARP_SIZE-1:0] mask);
        for(int i=0; i<WARP_SIZE; i++) if(mask[i]) return i;
        return 0;
    endfunction
    
    // Helper to count number of splits needed
    function automatic int count_splits(logic [WARP_SIZE-1:0] mask, logic [WARP_SIZE-1:0][31:0] addrs);
        logic [WARP_SIZE-1:0] remaining_mask;
        int split_count;
        int leader;
        
        remaining_mask = mask;
        split_count = 0;
        
        while (remaining_mask != 0) begin
            logic [WARP_SIZE-1:0] this_split_mask;
            leader = get_first_active_lane(remaining_mask);
            this_split_mask = '0;
            
            // Find all threads in same cache line as leader
            for (int i=0; i<WARP_SIZE; i++) begin
                if (remaining_mask[i] && (addrs[i][31:7] == addrs[leader][31:7])) begin
                    this_split_mask[i] = 1;
                end
            end
            
            remaining_mask = remaining_mask & ~this_split_mask;
            split_count++;
        end
        
        return split_count;
    endfunction
    
    // ========================================================================
    // Replay Arbiter (Round-Robin)
    // ========================================================================
    logic [WARP_ID_WIDTH-1:0] replay_rr_ptr;
    
    always_comb begin
        // Check which replays are valid and have TX IDs available
        for (int w=0; w<NUM_WARPS; w++) begin
            replay_valid[w] = replay_queue[w].valid && !tx_id_fifo_empty[w];
        end
        
        // Round-robin arbiter
        replay_grant_valid = 0;
        replay_granted_warp = replay_rr_ptr;
        
        for (int i=0; i<NUM_WARPS; i++) begin
            logic [WARP_ID_WIDTH-1:0] candidate;
            candidate = WARP_ID_WIDTH'( (32'(replay_rr_ptr) + 32'(i)) % 32'(NUM_WARPS) );
            if (replay_valid[candidate]) begin
                replay_grant_valid = 1;
                replay_granted_warp = candidate;
                break;
            end
        end
    end
    
    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            replay_rr_ptr <= 0;
        end else if (replay_grant_valid && mem_request_valid) begin
            // Advance round-robin pointer when replay issues
            replay_rr_ptr <= (replay_granted_warp + 1) % NUM_WARPS;
        end
    end
    
    // ========================================================================
    // Request Source Multiplexer (Replay vs New LSU)
    // ========================================================================
    always_comb begin
        // Priority: Replay > New LSU (finish in-progress splits first)
        if (replay_grant_valid) begin
            current_is_replay = 1;
            current_lsu_request.valid = 1;
            current_lsu_request.warp = replay_queue[replay_granted_warp].warp;
            current_lsu_request.rd = replay_queue[replay_granted_warp].rd;
            current_lsu_request.op = opcode_t'(replay_queue[replay_granted_warp].op);
            current_lsu_request.mask = replay_queue[replay_granted_warp].pending_mask;
            current_lsu_request.addresses = replay_queue[replay_granted_warp].addresses;
            current_lsu_request.store_data = replay_queue[replay_granted_warp].store_data;
        end else begin
            current_is_replay = 0;
            current_lsu_request = lsu_mem;
        end
    end
    
    // ========================================================================
    // Split Calculation
    // ========================================================================
    always_comb begin
        current_split_mask = '0;
        next_split_mask = '0;
        split_is_last = 1;
        split_leader = 0;
        mem_request_valid = 0;
        
        if (current_lsu_request.valid && (current_lsu_request.op == OP_LDR || current_lsu_request.op == OP_STR)) begin
            // 1. Find Leader
            split_leader = get_first_active_lane(current_lsu_request.mask);
            
            // 2. Determine Cache Line Agreement (128B aligned -> 7 LSBs ignored)
            for (int i=0; i<WARP_SIZE; i++) begin
                if (current_lsu_request.mask[i]) begin
                    if (current_lsu_request.addresses[i][31:7] == current_lsu_request.addresses[split_leader][31:7]) begin
                        current_split_mask[i] = 1;
                    end
                end
            end
            
            // 3. Calculate Remainder
            next_split_mask = current_lsu_request.mask & ~current_split_mask;
            split_is_last = (next_split_mask == 0);
            
            // 4. Request valid if TX ID available
            if (!tx_id_fifo_empty[current_lsu_request.warp]) begin
                mem_request_valid = 1;
            end
        end
    end
    
    // ========================================================================
    // Replay Queue Management
    // ========================================================================
    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            for (int w=0; w<NUM_WARPS; w++) begin
                replay_queue[w] <= '{valid:0, pending_mask:0, warp:0, rd:0, op:0, addresses:0, store_data:0};
            end
        end else begin
            // Update replay queue when requests are issued
            if (mem_request_valid) begin
                logic [WARP_ID_WIDTH-1:0] warp_idx;
                warp_idx = current_lsu_request.warp[WARP_ID_WIDTH-1:0];
                
                if (current_is_replay) begin
                    // Replay entry: update or clear
                    if (split_is_last) begin
                        replay_queue[warp_idx].valid <= 0;
                    end else begin
                        replay_queue[warp_idx].pending_mask <= next_split_mask;
                    end
                end else begin
                    // New LSU request: create replay if needed
                    if (!split_is_last) begin
                        replay_queue[warp_idx].valid <= 1;
                        replay_queue[warp_idx].pending_mask <= next_split_mask;
                        replay_queue[warp_idx].warp <= current_lsu_request.warp;
                        replay_queue[warp_idx].rd <= current_lsu_request.rd;
                        replay_queue[warp_idx].op <= current_lsu_request.op;
                        replay_queue[warp_idx].addresses <= current_lsu_request.addresses;
                        replay_queue[warp_idx].store_data <= current_lsu_request.store_data;
                    end
                end
            end
        end
    end

    // Shared Memory Signals
    logic shared_req_valid;
    logic shared_we;
    logic [WARP_SIZE-1:0] shared_req_mask;
    logic [WARP_SIZE-1:0][31:0] shared_rdata;

    // Shared Memory Pipeline Register (for 1-cycle latency)
    typedef struct packed {
        logic valid;
        logic [WARP_ID_WIDTH-1:0] warp;
        logic [REG_ADDR_WIDTH-1:0] rd;
        logic [WARP_SIZE-1:0] mask;
    } shared_wb_req_t;
    shared_wb_req_t shared_wb_req_q;

    typedef struct packed {
        logic valid;
        logic [WARP_ID_WIDTH-1:0] warp;
        logic [REG_ADDR_WIDTH-1:0] rd;
        logic [WARP_SIZE-1:0] mask;
        logic [WARP_SIZE-1:0][31:0] data;
    } shared_wb_resp_t;
    shared_wb_resp_t shared_wb_resp_q;



    // Output Registers from Cache Read
    logic [1023:0] l1_rdata_latched;

    // Address Conversion Logic (Word Index -> Byte Address)
    logic [WARP_SIZE-1:0][31:0] mem_addr_bytes;
    
    // Mock Memory Integration
    logic mock_req_valid;
    logic mock_req_ready;
    logic mock_resp_valid;
    logic [1023:0] mock_rdata;
    logic [WARP_ID_WIDTH-1:0]    mock_resp_warp;
    
    // ----------------------------------------------------------------
    // Simplified Packers (Assumes Coalesced Access for MVP/Test)
    // ----------------------------------------------------------------
    logic [31:0]   mock_base_addr;
    logic [1023:0] mock_wdata;
    logic [31:0]   mock_wmask;
    
    always_comb begin
        // 1. Calculate Base Address (from Split Leader)
        // Uses the aligned address of the first active lane in this split
        mock_base_addr = current_lsu_request.addresses[split_leader] & 32'hFFFFFF80;
        
        // 2. Pack Data & Mask (using current_split_mask)
        mock_wdata = '0;
        mock_wmask = '0;
        
        for (int i=0; i<WARP_SIZE; i++) begin
            if (current_split_mask[i]) begin
                logic [4:0] idx; 
                // idx = (Addr % 128) / 4
                idx = current_lsu_request.addresses[i][6:2]; 
                mock_wdata[idx*32 +: 32] = current_lsu_request.store_data[i];
                mock_wmask[idx] = 1;
            end
        end
    end

    // Use coalescer_valid signal from FSM as request trigger
    
    // Transaction ID signals
    logic [15:0] mock_req_transaction_id;
    logic [15:0] mock_resp_transaction_id;

    // Instantiate Mock Memory
    mock_memory dut_memory (
        .clk(clk),
        .rst_n(rst_n),
        .req_valid(mock_req_valid),
        .req_warp_id(lsu_mem.warp), // Pass Warp ID from LSU Pipeline
        .req_transaction_id(mock_req_transaction_id),
        .req_we(lsu_mem.op == OP_STR),
        .req_addr(mock_base_addr),
        .req_wdata(mock_wdata),
        .req_mask(mock_wmask),
        .req_ready(mock_req_ready),
        
        .resp_valid(mock_resp_valid),
        .resp_warp_id(mock_resp_warp),
        .resp_transaction_id(mock_resp_transaction_id),
        .resp_rdata(mock_rdata)
    );

    // Generate unique Request ID for Shared Memory based on instruction flow
    logic [7:0] lsu_req_toggle;
    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) lsu_req_toggle <= 0;
        else if (lsu_pop) lsu_req_toggle <= lsu_req_toggle + 1;
    end

    // Shared Memory (16KB) with Bank Conflict Serialization
    logic shared_mem_busy;
    logic [7:0] shared_conflict_cycles;
    
    shared_memory #(
        .SIZE_BYTES(16384),
        .NUM_BANKS(WARP_SIZE),
        .CONFLICT_MODE(2)  // 0=ignore, 1=warn, 2=serialize 
    ) local_memory (
        .clk(clk),
        .rst_n(rst_n),
        .req_valid(shared_req_valid),
        .req_uid({lsu_mem.op, lsu_req_toggle}), // Standard Toggle (No Lookahead)
        .req_mask(shared_req_mask),
        .req_we(shared_we),
        .req_addr(lsu_mem.addresses),
        .req_wdata(lsu_mem.store_data),
        .resp_rdata(shared_rdata),
        .busy(shared_mem_busy),
        .stall_cpu(shared_mem_stall_cpu),
        .conflict_cycles(shared_conflict_cycles)
    );
    
    // Connect Back to FSM Signals
    
    // Non-Blocking Adaptation:
    // We do NOT stall. We assume `mock_memory` handles the request.
    // We map the response directly to the Async Writeback logic.
    
    // Map L1 response signals for WB Consumption
    assign l1_resp_valid = mock_resp_valid; 
    assign mem_busy      = 0; // Never blocking
    assign l1_resp_rdata = mock_rdata; 
    // Stall Pipeline during Initialization Phase
    assign fsm_stall = (cycle < MAX_PENDING_PER_WARP + 5); 

    //=========================================================================
    // PIPELINE STAGE: WB (Writeback) + Async Memory Response Handler
    //=========================================================================
    // - Writes ALU results to register file (synchronous path)
    // - Handles asynchronous memory responses via MSHR lookup
    // - Clears scoreboard bits when writes complete
    // - Reclaims transaction IDs back to free pool
    //=========================================================================

    // Transaction ID Allocation
    logic mem_launch;
    
    // Memory launch condition: valid request from replay arbiter or new LSU
    // CRITICAL: mem_request_valid already checks TX ID availability
    assign mem_launch = mem_request_valid;
    
    // Shared Memory Launch
    assign shared_req_valid = lsu_mem.valid && (lsu_mem.op == OP_LDS || lsu_mem.op == OP_STS);
    assign shared_we        = (lsu_mem.op == OP_STS);
    assign shared_req_mask  = lsu_mem.mask;

    // Logic to issue request to Mock Memory
    assign mock_req_valid = mem_launch;
    assign coalescer_valid = mock_req_valid; // Alias if needed

    // ------------------------------------------------------------------------
    // UNIFIED MSHR & FIFO DRIVER LOGIC
    // ------------------------------------------------------------------------
    
    // Alloc Pop Logic (Combinational)
    always_comb begin
        for(int w=0; w<NUM_WARPS; w++) begin
             alloc_pop[w] = 0;
             if (mem_launch && lsu_mem.warp == 5'(w)) begin
                 alloc_pop[w] = 1;
             end
        end
    end
    
    // ------------------------------------------------------------------------
    // PATH C: FPU Pipeline (Execution & WB Stage)
    // ------------------------------------------------------------------------
    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            fpu_wb <= '{valid:0, src:WB_FPU, warp:0, rd:0, mask:0, result:0, we:0, we_pred:0, last_split:1, default:0};
        end else begin
            if (!stall_fpu_wb) begin 
                fpu_wb <= '{valid:0, src:WB_FPU, warp:0, rd:0, mask:0, result:0, we:0, we_pred:0, last_split:1, default:0}; // Removed op
                
                // --- SQUASH HANDLING ---
                if (fpu_inst_exec.branch_tag != warp_branch_tag[fpu_inst_exec.warp]) begin
                     // SQUASHED: Generate Dummy WB to clear Scoreboard
                     fpu_wb.valid <= 1;
                     fpu_wb.src   <= WB_SQUASH; // Tag as Squash
                     fpu_wb.warp  <= fpu_inst_exec.warp;
                     fpu_wb.rd    <= fpu_inst_exec.rd;
                     fpu_wb.mask  <= '0; // No side effects
                     fpu_wb.we    <= 0;  // No Register Write
                end else if (fpu_valid_exec) begin
                    
                    fpu_wb.valid <= 1;
                    fpu_wb.src   <= WB_FPU; // Tag as FPU
                    fpu_wb.warp  <= fpu_inst_exec.warp;
                    fpu_wb.rd    <= fpu_inst_exec.rd;
                    fpu_wb.mask  <= exec_mask_fpu; 
                    fpu_wb.we <= 1; 

                    if (fpu_inst_exec.op >= OP_SFU_SIN && fpu_inst_exec.op <= OP_SFU_TANH) begin
                        fpu_wb.result <= sfu_out_32b;
                    end else if (fpu_inst_exec.op == OP_FFMA || fpu_inst_exec.op == OP_FADD || fpu_inst_exec.op == OP_FMUL) begin
                        fpu_wb.result <= fma_out;
                    end else begin
                        // FSUB, ITOF etc use standard FPU/ALU
                        fpu_wb.result <= fpu_out;
                    end
                end
            end else begin
                // STALL: Hold fpu_wb state, do NOT update from pipeline
                // This will backpressure fpu_pop
            end
        end
    end

    // ------------------------------------------------------------------------
    // ATOMIC MEMORY WRITEBACK ARBITRATION (Combinational Next-State)
    // ------------------------------------------------------------------------
    logic global_mem_wb_ready;
    logic [WARP_ID_WIDTH-1:0] g_warp;
    int g_slot;
    pending_load_t g_info;
    
    always_comb begin
        g_warp = mock_resp_warp;
        g_slot = 32'(mock_resp_transaction_id[SLOT_ID_WIDTH-1:0]);
        global_mem_wb_ready = l1_resp_valid && (mshr_count[g_warp] > 0) && mshr_valid[g_warp][g_slot] && 
                             (mshr_table[g_warp][g_slot].transaction_id == mock_resp_transaction_id);
        g_info = mshr_table[g_warp][g_slot];

        mem_resp_wb_next = '{valid:0, src:WB_MEM, default:0};
        stall_shared_mem_wb = 0;

        // Priority 1: Global Memory Response (highest latency, critical)
        if (global_mem_wb_ready && !g_info.is_store) begin
            mem_resp_wb_next.valid    = 1;
            mem_resp_wb_next.src      = WB_MEM;
            mem_resp_wb_next.we       = 1;
            mem_resp_wb_next.warp     = g_warp;
            mem_resp_wb_next.rd       = {2'b0, g_info.rd[REG_ADDR_WIDTH-1:0]};
            mem_resp_wb_next.mask     = g_info.mask;
            mem_resp_wb_next.last_split = g_info.last_split;
            mem_resp_wb_next.we_pred  = 0;
            for (int l=0; l<WARP_SIZE; l++) begin
                if (g_info.mask[l]) begin
                    logic [4:0] idx = g_info.addresses[l][6:2];
                    mem_resp_wb_next.result[l] = l1_resp_rdata[idx*32 +: 32];
                end else begin
                    mem_resp_wb_next.result[l] = 32'h0;
                end
            end
            
            // Backpressure: If Global occupies WB, stall Shared pipeline
            if (shared_wb_resp_q.valid) stall_shared_mem_wb = 1;
        end
        // Priority 2: Shared Memory Response (2-Stage Pipelined)
        else if (shared_wb_resp_q.valid) begin
            mem_resp_wb_next.valid    = 1;
            mem_resp_wb_next.src      = WB_MEM;
            mem_resp_wb_next.we       = 1;
            mem_resp_wb_next.warp     = shared_wb_resp_q.warp;
            mem_resp_wb_next.rd       = {2'b0, shared_wb_resp_q.rd};
            mem_resp_wb_next.mask     = shared_wb_resp_q.mask;
            mem_resp_wb_next.result   = shared_wb_resp_q.data; 
            mem_resp_wb_next.last_split = 1; // Shared Mem is atomic for now
            mem_resp_wb_next.we_pred  = 0;
        end
        // Priority 3: Shadow NOP (Squash)
        else if (lsu_mem.valid && lsu_mem.op == OP_NOP) begin
            mem_resp_wb_next.valid    = 1;
            mem_resp_wb_next.src      = WB_SQUASH;
            mem_resp_wb_next.we       = 0; // Scoreboard clear only, no register write
            mem_resp_wb_next.warp     = lsu_mem.warp;
            mem_resp_wb_next.rd       = lsu_mem.rd;
            mem_resp_wb_next.mask     = '0;
            mem_resp_wb_next.last_split = 1; // Always clear on squash
            mem_resp_wb_next.we_pred  = 0;
            mem_resp_wb_next.result   = '0;
        end
    end

    // Consumption logic for stallable LSU pipeline
    assign lsu_mem_consumed = (lsu_mem.valid && lsu_mem.op == OP_NOP && mem_resp_wb_next.src == WB_SQUASH) || // Squash consumed only if WB granted
                              (lsu_mem.valid && (lsu_mem.op == OP_LDS || lsu_mem.op == OP_STS) && !shared_mem_stall_cpu && mem_resp_wb_next.valid) || // Shared consumed if no stall
                              (!current_is_replay && mem_request_valid); // New global request consumed if issued

    // ------------------------------------------------------------------------
    // LSU/MEM EXECUTION STAGE (Sequential)
    // ------------------------------------------------------------------------
    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            for(int w=0; w<NUM_WARPS; w++) begin
                reclaim_push[w] <= 0;
                mshr_valid[w] <= '0;
                mshr_count[w] <= 0;
            end
            async_wb_en <= 0;
            mem_resp_wb <= '{valid:0, src:WB_SQUASH, default:0};
            shared_wb_req_q <= '{valid:0, default:0};
            shared_wb_resp_q <= '{valid:0, default:0};
        end else begin
            // Register the Atomic Writeback Packet
            mem_resp_wb <= mem_resp_wb_next;

            // Default: Clear pulse signals
            for(int w=0; w<NUM_WARPS; w++) reclaim_push[w] <= 0;
            async_wb_en <= 0;
            
            if (shared_req_valid && !shared_mem_stall_cpu) begin
                shared_wb_req_q.valid <= 1;
                shared_wb_req_q.warp  <= lsu_mem.warp;
                shared_wb_req_q.rd    <= REG_ADDR_WIDTH'(lsu_mem.rd);
                shared_wb_req_q.mask  <= lsu_mem.mask;
            end else if (!stall_shared_mem_wb) begin
                shared_wb_req_q.valid <= 0;
            end
            
            // STAGE 2: Capture Data (1 cycle later)
            if (!stall_shared_mem_wb) begin
                shared_wb_resp_q.valid <= shared_wb_req_q.valid;
                shared_wb_resp_q.warp  <= shared_wb_req_q.warp;
                shared_wb_resp_q.rd    <= shared_wb_req_q.rd;
                // Explicitly cast or assign full width
                shared_wb_resp_q.mask  <= shared_wb_req_q.mask;
                shared_wb_resp_q.data  <= shared_rdata; 
            end

            // Allocation Logic (State Update Only)
            if (mem_launch) begin
                pending_load_t info;
                info.rd        = current_lsu_request.rd;
                // Use the SPLIT mask, not the full mask
                info.mask      = current_split_mask;
                info.last_split = split_is_last;
                info.is_store  = (current_lsu_request.op == OP_STR);
                info.transaction_id = mock_req_transaction_id;
                info.addresses = current_lsu_request.addresses;

                mshr_table[current_lsu_request.warp[WARP_ID_WIDTH-1:0]][mock_req_transaction_id[SLOT_ID_WIDTH-1:0]] <= info;
                mshr_valid[current_lsu_request.warp[WARP_ID_WIDTH-1:0]][mock_req_transaction_id[SLOT_ID_WIDTH-1:0]] <= 1;
                
                $display("CORE [%0t] TX_ID ALLOC: Warp=%0d TxID=%0d Store=%b Mask=%h", 
                         $time, current_lsu_request.warp, mock_req_transaction_id, info.is_store, info.mask);
            end


        // -----------------------
        // RECLAMATION LOGIC (Priority 1)
        // -----------------------
            // Reclamation Logic (State updates only - data is handled by mem_resp_wb_next)
            if (global_mem_wb_ready) begin
                reclaim_data[g_warp] <= g_info.transaction_id;
                reclaim_push[g_warp] <= 1;
                mshr_valid[g_warp][g_slot] <= 0;
                
                if (!g_info.is_store) begin
                    async_wb_en   <= 1;
                    async_wb_warp <= g_warp;
                    async_wb_rd   <= g_info.rd;
                end
            end

        
        // -----------------------
        // MSHR COUNT UPDATE (Safe Merge)
        // -----------------------
        for (int w=0; w<NUM_WARPS; w++) begin
            int next_cnt;
            logic [WARP_ID_WIDTH-1:0] cur_w;
            cur_w = WARP_ID_WIDTH'(w);
            next_cnt = mshr_count[cur_w];
            
            // Increment if Allocating (Correctly identify the issued warp)
            // MUST NOT be gated by stall_pipeline because the launch to mock memory is NOT gated.
            if (mem_launch && current_lsu_request.warp == cur_w)
                next_cnt++;
                
            // Decrement if Reclaiming
            if (l1_resp_valid && mock_resp_warp == cur_w && mshr_count[cur_w] > 0) begin
                logic [SLOT_ID_WIDTH-1:0] q_idx;
                q_idx = mock_resp_transaction_id[SLOT_ID_WIDTH-1:0];
                if (mshr_valid[cur_w][q_idx] && mshr_table[cur_w][q_idx].transaction_id == mock_resp_transaction_id)
                    next_cnt--;
            end
                
            mshr_count[cur_w] <= next_cnt;
        end
        
        // -----------------------
        // PIPELINE WRITEBACK (Priority 2)
        // -----------------------
        if (mem_wb.valid && mem_wb.we) begin
            // Sync writeback logic is now handled by oc_wb[0] assignment (combinational or driven by OC)
            // Removed redundant direct GPR writes
        end
        end
    end
    
    // Drive transaction ID to mock_memory (peek at what we're about to pop)
    // This is safe because we only peek when mem_launch is true (same condition as pop)
    assign mock_req_transaction_id = (mem_launch) ?
                                      tx_id_fifo_dout[lsu_mem.warp[WARP_ID_WIDTH-1:0]] :  // Peek at front of LSU warp's FIFO
                                      16'h0;

    // Simulation Control & Initialization

    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            cycle <= 0;
            done  <= 0;
            done_prev <= 0;
            done_prev <= 0;
            barrier_mask       <= 0;
            barrier_expected   <= 0; // Initialize to 0, latch active warps below
            barrier_epoch      <= 0;
            barrier_seen_epoch <= 0;
            barrier_active     <= 0;
            barrier_initialized <= 0;
            
            // Initialize MSHR tables
            // MSHR Init moved to Unified Driver
            
            // Clear Init Signals
            for (int w=0; w<NUM_WARPS; w++) begin
                init_push[w] <= 0;
            end
            
            for (int w=0; w<NUM_WARPS; w++) begin
                // All architectural state is now managed and reset in the 
                // relevant pipeline stage blocks (Scheduler, ID) to avoid multiple drivers.
                // init_push and other memory-related signals are still reset here.
                init_push[w] <= 0;
            end
        end else begin
            // Populate TX ID FIFOs over first MAX_PENDING_PER_WARP cycles
            if (cycle < MAX_PENDING_PER_WARP) begin
                for (int w=0; w<NUM_WARPS; w++) begin
                    logic [TX_ID_WIDTH-1:0] tx_id;
                    tx_id = '0;
                    tx_id[SM_ID_OFFSET +: 4] = SM_ID[3:0];
                    tx_id[WARP_ID_OFFSET +: WARP_ID_WIDTH] = w[WARP_ID_WIDTH-1:0];
                    tx_id[0 +: SLOT_ID_WIDTH] = cycle[SLOT_ID_WIDTH-1:0];
                    
                    init_data[w] <= tx_id;
                    init_push[w] <= 1;
                end
            end else if (cycle == MAX_PENDING_PER_WARP) begin
                // Clear Push after Init
                for (int w=0; w<NUM_WARPS; w++) begin
                    init_push[w] <= 0;
                end
                $display("INIT: Populated TX ID FIFOs for %0d warps with %0d IDs each", 
                         NUM_WARPS, MAX_PENDING_PER_WARP);
            end
            
            cycle <= cycle + 1;
            
            init_phase <= (cycle < MAX_PENDING_PER_WARP + 2);
            done       <= done_next;
            if (done && !done_prev) $display("CORE [%0t] ALL WARPS EXITED", $time);
            done_prev  <= done;

            // BREAK COMBINATIONAL LOOPS
            // 1. Register Scoreboard Clears
            reg_clear_q <= reg_clear_this_cycle;

            // 2. Register Writeback Port Control (Stability for OC)
            for (int k=0; k<2; k++) begin
                oc_wb_valid_q[k]   <= oc_wb_valid[k];
                oc_wb_warp_q[k]    <= oc_wb_warp[k];
                oc_wb_rd_q[k]      <= oc_wb_rd[k];
                oc_wb_mask_q[k]    <= oc_wb_mask[k];
                oc_wb_result_q[k]  <= oc_wb_data[k];
                oc_wb_we_q[k]      <= 1'b1; // Default - data carries actual mask
                // Special case for we_pred if needed, currently results carry mask
            end
        end
    end

    // Stable done calculation
    always_comb begin
        done_next = 1;
        for (int w=0; w<NUM_WARPS; w++) begin
            if (warp_state[w] != W_EXIT && warp_state[w] != W_IDLE) begin
                done_next = 0;
            end
        end
    end

    // DEDICATED EX -> IF BRANCH REGISTER BLOCK
    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            branch_taken_q  <= 0;
            branch_warp_q   <= 0;
            branch_target_q <= 0;
        end else begin
            branch_taken_q  <= cur_branch_taken;
            branch_warp_q   <= cur_branch_warp;
            branch_target_q <= cur_branch_target;
        end
    end
    // COMPREHENSIVE ASSERTION BLOCK (Transaction ID Allocator)

    // Validates free list integrity and catches allocation/reclamation bugs
    // All complex assertions with variable declarations are here to avoid syntax issues

    
    always_ff @(posedge clk) begin
        if (rst_n) begin
            // PERIODIC INVARIANT CHECKS (Every Cycle)
            for (int w = 0; w < NUM_WARPS; w++) begin
                if (cycle > MAX_PENDING_PER_WARP + 10) begin
                    int total_ids;
                    total_ids = int'(tx_id_fifo_count[w]) + mshr_count[w] + int'(reclaim_push[w]) - int'(alloc_pop[w]);
                    
                    if (total_ids != MAX_PENDING_PER_WARP) begin
                        // Relaxed: Just print warning instead of stop
                        $display("CORE [%0t] INVARIANT WARNING: Warp %0d has %0d(fifo) + %0d(mshr) + %0d(rec) - %0d(alloc) = %0d (expected %0d)",
                               $time, w, tx_id_fifo_count[w], mshr_count[w], reclaim_push[w], alloc_pop[w],
                               total_ids, MAX_PENDING_PER_WARP);
                    end
                end
                
                // INVARIANT 2: All free list IDs belong to this SM and warp's partition
                // (Cannot peek into FIFO for all elements easily - skipping)
                
                // INVARIANT 3: Free list size never exceeds MAX_PENDING_PER_WARP
                assert (tx_id_fifo_count[w] <= MAX_PENDING_PER_WARP) else
                    $fatal(1, "CORE [%0t] FREE LIST OVERFLOW: Warp %0d has %0d IDs (max %0d)",
                           $time, w, tx_id_fifo_count[w], MAX_PENDING_PER_WARP);
            end
        end
    end

    // Helper Functions
    function automatic [31:0] count_leading_zeros(input [31:0] in);
        for (int i=31; i>=0; i--) begin
            if (in[i]) return 31-i;
        end
        return 32;
    endfunction

    function automatic [31:0] double_to_float(input [63:0] d);
        logic sign;
        logic [10:0] exp64;
        logic [51:0] mant64;
        logic [7:0] exp32;
        logic [22:0] mant32;

        sign = d[63];
        exp64 = d[62:52];
        mant64 = d[51:0];

        if (exp64 == 0) return 32'b0; // Zero
        // Simplified conversion: doesn't handle Inf/NaN/Denorm perfectly but works for normal integers
        
        exp32 = 8'(exp64 - 11'd1023 + 11'd127);
        mant32 = mant64[51:29]; 

        return {sign, exp32, mant32};
    endfunction

    // ASSERTION: Double WB Owner Check
    always_ff @(posedge clk) begin
        if (rst_n) begin
            // Check if multiple sources are trying to WB to the same warp/reg
            // We ignore Rd 0 as it is often a dummy destination for squashed/non-writing ops
            // Must check WE (Write Enable) to actual data conflicts (Squashed insts have valid=1 but we=0)
            if (alu_wb.valid && alu_wb.we && mem_resp_wb.valid && mem_resp_wb.we && alu_wb.warp == mem_resp_wb.warp && alu_wb.rd == mem_resp_wb.rd && alu_wb.rd != 0)
                    $fatal(1, "CORE [%0t] DOUBLE WB OWNER: Warp %0d Rd %0d (ALU vs MEM)", $time, alu_wb.warp, alu_wb.rd);
            if (fpu_wb.valid && fpu_wb.we && mem_resp_wb.valid && mem_resp_wb.we && fpu_wb.warp == mem_resp_wb.warp && fpu_wb.rd == mem_resp_wb.rd && fpu_wb.rd != 0)
                    $fatal(1, "CORE [%0t] DOUBLE WB OWNER: Warp %0d Rd %0d (FPU vs MEM)", $time, fpu_wb.warp, fpu_wb.rd);
        end
    end

    // CENTRALIZED WARP STATE DRIVER
    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            for (int w=0; w<NUM_WARPS; w++) begin
                warp_state[w] <= W_IDLE;
            end
        end else begin
            for (int w=0; w<NUM_WARPS; w++) begin
                warp_state[w] <= warp_state_next[w];
            end
        end
    end

    // WARP STATE NEXT-STATE LOGIC
    always_comb begin
        for (int w=0; w<NUM_WARPS; w++) begin
            warp_state_next[w] = warp_state[w];
            
            // Priority 1: Exit Request
            if (state_req_exit[w]) begin
                warp_state_next[w] = W_EXIT;
            end
            // Priority 2: Ready Request (Barrier Release)
            else if (state_req_ready[w]) begin
                warp_state_next[w] = W_READY;
            end
            // Priority 3: Barrier Request (Arrive at Barrier)
            else if (state_req_barrier[w]) begin
                warp_state_next[w] = W_BARRIER;
            end
        end
    end

    // STUBS FOR DISTRIBUTED STATE REQUESTS (Combinational)
    always_comb begin
        state_req_exit    = '0;
        state_req_barrier = '0;
        state_req_ready   = '0;

        // ALU EX Stage: EXIT (Waits for MSHR Drain for Consistency)
        if (alu_valid_exec && alu_can_commit && (alu_inst_exec.branch_tag == warp_branch_tag[alu_inst_exec.warp])) begin
            if (alu_inst_exec.op == OP_EXIT) begin
                // Ensure all pending memory transactions (Shared/Global) are complete
                // AND written back (cover pipeline latency MSHR -> WB)
                logic pipeline_busy;
                pipeline_busy = (mshr_count[alu_inst_exec.warp] != 0) ||
                                (lsu_valid_exec && lsu_inst_exec.warp == alu_inst_exec.warp) || // Sibling LSU op
                                (lsu_mem.valid && lsu_mem.warp == alu_inst_exec.warp) ||        // MEM stage
                                (shared_wb_resp_q.valid && shared_wb_resp_q.warp == alu_inst_exec.warp) || // Shared WB
                                (mem_resp_wb.valid && mem_resp_wb.warp == alu_inst_exec.warp) || // Global WB
                                (oc_wb_valid_q[0] && oc_wb_warp_q[0] == alu_inst_exec.warp) ||   // RF Write Port 0
                                (oc_wb_valid_q[1] && oc_wb_warp_q[1] == alu_inst_exec.warp);     // RF Write Port 1

                if (!pipeline_busy) begin
                    state_req_exit[alu_inst_exec.warp] = 1;
                end
            end
        end

        // ALU EX Stage: BAR Arrival (Waits for MSHR Drain for Consistency)
        if (alu_valid_exec && alu_can_commit && (alu_inst_exec.branch_tag == warp_branch_tag[alu_inst_exec.warp])) begin
            if (alu_inst_exec.op == OP_BAR) begin
                // Memory Consistency: Ensure all previous loads have retired
                if (mshr_count[alu_inst_exec.warp] == 0) begin
                    if (barrier_seen_epoch[alu_inst_exec.warp] != barrier_epoch) begin
                        state_req_barrier[alu_inst_exec.warp] = 1;
                    end
                end
            end
        end

        // Barrier Logic: RELEASE
        if (barrier_initialized && 
            ((barrier_mask | (1 << alu_inst_exec.warp)) & barrier_expected) == barrier_expected && barrier_expected != 0) begin
            if (alu_inst_exec.op == OP_BAR) begin
                for (int i = 0; i < NUM_WARPS; i++) begin
                    if (barrier_expected[i] && warp_state[i] == W_BARRIER)
                        state_req_ready[i] = 1;
                end
                state_req_ready[alu_inst_exec.warp] = 1;
            end
        end
    end

    // Warp 7 diagnostic block
    always_ff @(posedge clk) begin
        static int cycle_diag = 0;
        cycle_diag++;
        if (cycle_diag % 100 == 0) begin
            $display("CORE [%0t] WARP7_DIAG: PC=%h State=%s SB=%b PredSB=%b MSHR=%d", 
                     $time, warp_pc[7], warp_state[7].name(), warp_reg_writes[7], warp_pred_writes[7], mshr_count[7]);
        end
    end
endmodule
